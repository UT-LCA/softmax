module logunit (a, z, status);
	
	input [31:0] a;
	output reg [31:0] z;
	output [7:0] status;

	wire [28: 0] fx;
	wire [31: 0] fxout1;
	wire [31: 0] fxout2;
	wire [31:0] temp;	

	fptofixed_para fptofx(.fp(a),.fx(fx));
	LUT1 lut1 (.addr(fx[27:23]),.log(fxout1)); 
	LUT2 lut2 (.addr(fx[22:11]),.log(fxout2));  
	DW01_add #(32) addsub1 (.A(fxout1),.B(fxout2),.CI(1'b0),.SUM(temp),.CO());

always @(temp)
begin
	if (fx[28] == 1) z <= 32'h80000001;
	else z <= temp;
end
endmodule

module fptofixed_para (
	fp,
	fx
	);
	
	

	input [31:0] fp; // Half Precision fp
	output [28:0] fx;  
	
	wire [31:0] dec;
	wire [5:0] enc;


	wire [30:0] temp;
	//wire grt;
	wire [30:0] temp2;
	reg [31:0] temp3;

	assign temp = fp[30:0];
	assign fx = {enc,temp3[30:8]};

always @(temp2)
begin
	if (dec[31:0] == 0)
		begin
			temp3 <= 31'h00000000;		
		end

	else 
		begin
			temp3 <= temp2;
		end
end	

DW_lzd #(32) lzd (.a(fp),.enc(enc),.dec(dec));
DW01_ash #(31,6) ash( .A(temp[30:0]), .DATA_TC(1'b0), .SH(enc), .SH_TC(1'b0), .B(temp2));
//DW01_addsub #(32) addsub1 (.A(fp),.B(32'h00000001),.CI(1'b0),.ADD_SUB(1'b1),.SUM(temp),.CO());
endmodule

module LUT1(addr, log);
    input [4:0] addr;
    output reg [31:0] log;

    always @(addr) begin
        case (addr)
			5'b0 		: log = 32'b00000000000010100110010110101111;
			5'b1 		: log = 32'b00000000000010011011010000111101;
			5'b10 		: log = 32'b00000000000010010000001011001011;
			5'b11 		: log = 32'b00000000000010000101000101011001;
			5'b100 		: log = 32'b00000000000001111001111111100111;
			5'b101 		: log = 32'b00000000000001101110111001110100;
			5'b110 		: log = 32'b00000000000001100011110100000010;
			5'b111 		: log = 32'b00000000000001011000101110010000;
			5'b1000 		: log = 32'b00000000000001001101101000011110;
			5'b1001 		: log = 32'b00000000000001000010100010101100;
			5'b1010 		: log = 32'b00000000000000110111011100111010;
			5'b1011 		: log = 32'b00000000000000101100010111001000;
			5'b1100 		: log = 32'b00000000000000100001010001010110;
			5'b1101 		: log = 32'b00000000000000010110001011100100;
			5'b1110 		: log = 32'b00000000000000001011000101110010;
			5'b1111 		: log = 32'b00000000000000000000000000000000;
			5'b10000 		: log = 32'b11111111111111111011000101110010;
			5'b10001 		: log = 32'b11111111111111110110001011100100;
			5'b10010 		: log = 32'b11111111111111100001010001010110;
			5'b10011 		: log = 32'b11111111111111101100010111001000;
			5'b10100 		: log = 32'b11111111111111110111011100111010;
			5'b10101 		: log = 32'b11111111111111000010100010101100;
			5'b10110 		: log = 32'b11111111111111001101101000011110;
			5'b10111 		: log = 32'b11111111111111011000101110010000;
			5'b11000 		: log = 32'b11111111111111100011110100000010;
			5'b11001 		: log = 32'b11111111111111101110111001110100;
			5'b11010 		: log = 32'b11111111111111111001111111100111;
			5'b11011 		: log = 32'b11111111111110000101000101011001;
			5'b11100 		: log = 32'b11111111111110010000001011001011;
			5'b11101 		: log = 32'b11111111111110011011010000111101;
			5'b11110 		: log = 32'b11111111111110100110010110101111;
			5'b11111 		: log = 32'b11111111111110110001011100100001;
        endcase
    end
endmodule

module LUT2(addr, log);
    input [11:0] addr;
    output reg [31:0] log;

    always @(addr) begin
        case (addr)
			12'b0 		: log = 32'b00000000000000000000000000000000;
			12'b1 		: log = 32'b00000000000000000000000000001111;
			12'b10 		: log = 32'b00000000000000000000000000011111;
			12'b11 		: log = 32'b00000000000000000000000000101111;
			12'b100 		: log = 32'b00000000000000000000000000111111;
			12'b101 		: log = 32'b00000000000000000000000001001111;
			12'b110 		: log = 32'b00000000000000000000000001011111;
			12'b111 		: log = 32'b00000000000000000000000001101111;
			12'b1000 		: log = 32'b00000000000000000000000001111111;
			12'b1001 		: log = 32'b00000000000000000000000010001111;
			12'b1010 		: log = 32'b00000000000000000000000010011111;
			12'b1011 		: log = 32'b00000000000000000000000010101111;
			12'b1100 		: log = 32'b00000000000000000000000010111111;
			12'b1101 		: log = 32'b00000000000000000000000011001111;
			12'b1110 		: log = 32'b00000000000000000000000011011111;
			12'b1111 		: log = 32'b00000000000000000000000011101111;
			12'b10000 		: log = 32'b00000000000000000000000011111111;
			12'b10001 		: log = 32'b00000000000000000000000100001111;
			12'b10010 		: log = 32'b00000000000000000000000100011111;
			12'b10011 		: log = 32'b00000000000000000000000100101111;
			12'b10100 		: log = 32'b00000000000000000000000100111111;
			12'b10101 		: log = 32'b00000000000000000000000101001111;
			12'b10110 		: log = 32'b00000000000000000000000101011111;
			12'b10111 		: log = 32'b00000000000000000000000101101110;
			12'b11000 		: log = 32'b00000000000000000000000101111110;
			12'b11001 		: log = 32'b00000000000000000000000110001110;
			12'b11010 		: log = 32'b00000000000000000000000110011110;
			12'b11011 		: log = 32'b00000000000000000000000110101110;
			12'b11100 		: log = 32'b00000000000000000000000110111110;
			12'b11101 		: log = 32'b00000000000000000000000111001110;
			12'b11110 		: log = 32'b00000000000000000000000111011110;
			12'b11111 		: log = 32'b00000000000000000000000111101110;
			12'b100000 		: log = 32'b00000000000000000000000111111110;
			12'b100001 		: log = 32'b00000000000000000000001000001101;
			12'b100010 		: log = 32'b00000000000000000000001000011101;
			12'b100011 		: log = 32'b00000000000000000000001000101101;
			12'b100100 		: log = 32'b00000000000000000000001000111101;
			12'b100101 		: log = 32'b00000000000000000000001001001101;
			12'b100110 		: log = 32'b00000000000000000000001001011101;
			12'b100111 		: log = 32'b00000000000000000000001001101101;
			12'b101000 		: log = 32'b00000000000000000000001001111100;
			12'b101001 		: log = 32'b00000000000000000000001010001100;
			12'b101010 		: log = 32'b00000000000000000000001010011100;
			12'b101011 		: log = 32'b00000000000000000000001010101100;
			12'b101100 		: log = 32'b00000000000000000000001010111100;
			12'b101101 		: log = 32'b00000000000000000000001011001100;
			12'b101110 		: log = 32'b00000000000000000000001011011011;
			12'b101111 		: log = 32'b00000000000000000000001011101011;
			12'b110000 		: log = 32'b00000000000000000000001011111011;
			12'b110001 		: log = 32'b00000000000000000000001100001011;
			12'b110010 		: log = 32'b00000000000000000000001100011011;
			12'b110011 		: log = 32'b00000000000000000000001100101010;
			12'b110100 		: log = 32'b00000000000000000000001100111010;
			12'b110101 		: log = 32'b00000000000000000000001101001010;
			12'b110110 		: log = 32'b00000000000000000000001101011010;
			12'b110111 		: log = 32'b00000000000000000000001101101010;
			12'b111000 		: log = 32'b00000000000000000000001101111001;
			12'b111001 		: log = 32'b00000000000000000000001110001001;
			12'b111010 		: log = 32'b00000000000000000000001110011001;
			12'b111011 		: log = 32'b00000000000000000000001110101001;
			12'b111100 		: log = 32'b00000000000000000000001110111001;
			12'b111101 		: log = 32'b00000000000000000000001111001000;
			12'b111110 		: log = 32'b00000000000000000000001111011000;
			12'b111111 		: log = 32'b00000000000000000000001111101000;
			12'b1000000 		: log = 32'b00000000000000000000001111111000;
			12'b1000001 		: log = 32'b00000000000000000000010000000111;
			12'b1000010 		: log = 32'b00000000000000000000010000010111;
			12'b1000011 		: log = 32'b00000000000000000000010000100111;
			12'b1000100 		: log = 32'b00000000000000000000010000110111;
			12'b1000101 		: log = 32'b00000000000000000000010001000110;
			12'b1000110 		: log = 32'b00000000000000000000010001010110;
			12'b1000111 		: log = 32'b00000000000000000000010001100110;
			12'b1001000 		: log = 32'b00000000000000000000010001110101;
			12'b1001001 		: log = 32'b00000000000000000000010010000101;
			12'b1001010 		: log = 32'b00000000000000000000010010010101;
			12'b1001011 		: log = 32'b00000000000000000000010010100101;
			12'b1001100 		: log = 32'b00000000000000000000010010110100;
			12'b1001101 		: log = 32'b00000000000000000000010011000100;
			12'b1001110 		: log = 32'b00000000000000000000010011010100;
			12'b1001111 		: log = 32'b00000000000000000000010011100011;
			12'b1010000 		: log = 32'b00000000000000000000010011110011;
			12'b1010001 		: log = 32'b00000000000000000000010100000011;
			12'b1010010 		: log = 32'b00000000000000000000010100010011;
			12'b1010011 		: log = 32'b00000000000000000000010100100010;
			12'b1010100 		: log = 32'b00000000000000000000010100110010;
			12'b1010101 		: log = 32'b00000000000000000000010101000010;
			12'b1010110 		: log = 32'b00000000000000000000010101010001;
			12'b1010111 		: log = 32'b00000000000000000000010101100001;
			12'b1011000 		: log = 32'b00000000000000000000010101110001;
			12'b1011001 		: log = 32'b00000000000000000000010110000000;
			12'b1011010 		: log = 32'b00000000000000000000010110010000;
			12'b1011011 		: log = 32'b00000000000000000000010110100000;
			12'b1011100 		: log = 32'b00000000000000000000010110101111;
			12'b1011101 		: log = 32'b00000000000000000000010110111111;
			12'b1011110 		: log = 32'b00000000000000000000010111001111;
			12'b1011111 		: log = 32'b00000000000000000000010111011110;
			12'b1100000 		: log = 32'b00000000000000000000010111101110;
			12'b1100001 		: log = 32'b00000000000000000000010111111101;
			12'b1100010 		: log = 32'b00000000000000000000011000001101;
			12'b1100011 		: log = 32'b00000000000000000000011000011101;
			12'b1100100 		: log = 32'b00000000000000000000011000101100;
			12'b1100101 		: log = 32'b00000000000000000000011000111100;
			12'b1100110 		: log = 32'b00000000000000000000011001001100;
			12'b1100111 		: log = 32'b00000000000000000000011001011011;
			12'b1101000 		: log = 32'b00000000000000000000011001101011;
			12'b1101001 		: log = 32'b00000000000000000000011001111010;
			12'b1101010 		: log = 32'b00000000000000000000011010001010;
			12'b1101011 		: log = 32'b00000000000000000000011010011010;
			12'b1101100 		: log = 32'b00000000000000000000011010101001;
			12'b1101101 		: log = 32'b00000000000000000000011010111001;
			12'b1101110 		: log = 32'b00000000000000000000011011001000;
			12'b1101111 		: log = 32'b00000000000000000000011011011000;
			12'b1110000 		: log = 32'b00000000000000000000011011100111;
			12'b1110001 		: log = 32'b00000000000000000000011011110111;
			12'b1110010 		: log = 32'b00000000000000000000011100000111;
			12'b1110011 		: log = 32'b00000000000000000000011100010110;
			12'b1110100 		: log = 32'b00000000000000000000011100100110;
			12'b1110101 		: log = 32'b00000000000000000000011100110101;
			12'b1110110 		: log = 32'b00000000000000000000011101000101;
			12'b1110111 		: log = 32'b00000000000000000000011101010100;
			12'b1111000 		: log = 32'b00000000000000000000011101100100;
			12'b1111001 		: log = 32'b00000000000000000000011101110011;
			12'b1111010 		: log = 32'b00000000000000000000011110000011;
			12'b1111011 		: log = 32'b00000000000000000000011110010011;
			12'b1111100 		: log = 32'b00000000000000000000011110100010;
			12'b1111101 		: log = 32'b00000000000000000000011110110010;
			12'b1111110 		: log = 32'b00000000000000000000011111000001;
			12'b1111111 		: log = 32'b00000000000000000000011111010001;
			12'b10000000 		: log = 32'b00000000000000000000011111100000;
			12'b10000001 		: log = 32'b00000000000000000000011111110000;
			12'b10000010 		: log = 32'b00000000000000000000011111111111;
			12'b10000011 		: log = 32'b00000000000000000000100000001111;
			12'b10000100 		: log = 32'b00000000000000000000100000011110;
			12'b10000101 		: log = 32'b00000000000000000000100000101110;
			12'b10000110 		: log = 32'b00000000000000000000100000111101;
			12'b10000111 		: log = 32'b00000000000000000000100001001101;
			12'b10001000 		: log = 32'b00000000000000000000100001011100;
			12'b10001001 		: log = 32'b00000000000000000000100001101100;
			12'b10001010 		: log = 32'b00000000000000000000100001111011;
			12'b10001011 		: log = 32'b00000000000000000000100010001011;
			12'b10001100 		: log = 32'b00000000000000000000100010011010;
			12'b10001101 		: log = 32'b00000000000000000000100010101010;
			12'b10001110 		: log = 32'b00000000000000000000100010111001;
			12'b10001111 		: log = 32'b00000000000000000000100011001000;
			12'b10010000 		: log = 32'b00000000000000000000100011011000;
			12'b10010001 		: log = 32'b00000000000000000000100011100111;
			12'b10010010 		: log = 32'b00000000000000000000100011110111;
			12'b10010011 		: log = 32'b00000000000000000000100100000110;
			12'b10010100 		: log = 32'b00000000000000000000100100010110;
			12'b10010101 		: log = 32'b00000000000000000000100100100101;
			12'b10010110 		: log = 32'b00000000000000000000100100110101;
			12'b10010111 		: log = 32'b00000000000000000000100101000100;
			12'b10011000 		: log = 32'b00000000000000000000100101010011;
			12'b10011001 		: log = 32'b00000000000000000000100101100011;
			12'b10011010 		: log = 32'b00000000000000000000100101110010;
			12'b10011011 		: log = 32'b00000000000000000000100110000010;
			12'b10011100 		: log = 32'b00000000000000000000100110010001;
			12'b10011101 		: log = 32'b00000000000000000000100110100001;
			12'b10011110 		: log = 32'b00000000000000000000100110110000;
			12'b10011111 		: log = 32'b00000000000000000000100110111111;
			12'b10100000 		: log = 32'b00000000000000000000100111001111;
			12'b10100001 		: log = 32'b00000000000000000000100111011110;
			12'b10100010 		: log = 32'b00000000000000000000100111101110;
			12'b10100011 		: log = 32'b00000000000000000000100111111101;
			12'b10100100 		: log = 32'b00000000000000000000101000001100;
			12'b10100101 		: log = 32'b00000000000000000000101000011100;
			12'b10100110 		: log = 32'b00000000000000000000101000101011;
			12'b10100111 		: log = 32'b00000000000000000000101000111010;
			12'b10101000 		: log = 32'b00000000000000000000101001001010;
			12'b10101001 		: log = 32'b00000000000000000000101001011001;
			12'b10101010 		: log = 32'b00000000000000000000101001101001;
			12'b10101011 		: log = 32'b00000000000000000000101001111000;
			12'b10101100 		: log = 32'b00000000000000000000101010000111;
			12'b10101101 		: log = 32'b00000000000000000000101010010111;
			12'b10101110 		: log = 32'b00000000000000000000101010100110;
			12'b10101111 		: log = 32'b00000000000000000000101010110101;
			12'b10110000 		: log = 32'b00000000000000000000101011000101;
			12'b10110001 		: log = 32'b00000000000000000000101011010100;
			12'b10110010 		: log = 32'b00000000000000000000101011100011;
			12'b10110011 		: log = 32'b00000000000000000000101011110011;
			12'b10110100 		: log = 32'b00000000000000000000101100000010;
			12'b10110101 		: log = 32'b00000000000000000000101100010001;
			12'b10110110 		: log = 32'b00000000000000000000101100100001;
			12'b10110111 		: log = 32'b00000000000000000000101100110000;
			12'b10111000 		: log = 32'b00000000000000000000101100111111;
			12'b10111001 		: log = 32'b00000000000000000000101101001111;
			12'b10111010 		: log = 32'b00000000000000000000101101011110;
			12'b10111011 		: log = 32'b00000000000000000000101101101101;
			12'b10111100 		: log = 32'b00000000000000000000101101111101;
			12'b10111101 		: log = 32'b00000000000000000000101110001100;
			12'b10111110 		: log = 32'b00000000000000000000101110011011;
			12'b10111111 		: log = 32'b00000000000000000000101110101010;
			12'b11000000 		: log = 32'b00000000000000000000101110111010;
			12'b11000001 		: log = 32'b00000000000000000000101111001001;
			12'b11000010 		: log = 32'b00000000000000000000101111011000;
			12'b11000011 		: log = 32'b00000000000000000000101111101000;
			12'b11000100 		: log = 32'b00000000000000000000101111110111;
			12'b11000101 		: log = 32'b00000000000000000000110000000110;
			12'b11000110 		: log = 32'b00000000000000000000110000010101;
			12'b11000111 		: log = 32'b00000000000000000000110000100101;
			12'b11001000 		: log = 32'b00000000000000000000110000110100;
			12'b11001001 		: log = 32'b00000000000000000000110001000011;
			12'b11001010 		: log = 32'b00000000000000000000110001010010;
			12'b11001011 		: log = 32'b00000000000000000000110001100010;
			12'b11001100 		: log = 32'b00000000000000000000110001110001;
			12'b11001101 		: log = 32'b00000000000000000000110010000000;
			12'b11001110 		: log = 32'b00000000000000000000110010001111;
			12'b11001111 		: log = 32'b00000000000000000000110010011111;
			12'b11010000 		: log = 32'b00000000000000000000110010101110;
			12'b11010001 		: log = 32'b00000000000000000000110010111101;
			12'b11010010 		: log = 32'b00000000000000000000110011001100;
			12'b11010011 		: log = 32'b00000000000000000000110011011011;
			12'b11010100 		: log = 32'b00000000000000000000110011101011;
			12'b11010101 		: log = 32'b00000000000000000000110011111010;
			12'b11010110 		: log = 32'b00000000000000000000110100001001;
			12'b11010111 		: log = 32'b00000000000000000000110100011000;
			12'b11011000 		: log = 32'b00000000000000000000110100100111;
			12'b11011001 		: log = 32'b00000000000000000000110100110111;
			12'b11011010 		: log = 32'b00000000000000000000110101000110;
			12'b11011011 		: log = 32'b00000000000000000000110101010101;
			12'b11011100 		: log = 32'b00000000000000000000110101100100;
			12'b11011101 		: log = 32'b00000000000000000000110101110011;
			12'b11011110 		: log = 32'b00000000000000000000110110000011;
			12'b11011111 		: log = 32'b00000000000000000000110110010010;
			12'b11100000 		: log = 32'b00000000000000000000110110100001;
			12'b11100001 		: log = 32'b00000000000000000000110110110000;
			12'b11100010 		: log = 32'b00000000000000000000110110111111;
			12'b11100011 		: log = 32'b00000000000000000000110111001110;
			12'b11100100 		: log = 32'b00000000000000000000110111011110;
			12'b11100101 		: log = 32'b00000000000000000000110111101101;
			12'b11100110 		: log = 32'b00000000000000000000110111111100;
			12'b11100111 		: log = 32'b00000000000000000000111000001011;
			12'b11101000 		: log = 32'b00000000000000000000111000011010;
			12'b11101001 		: log = 32'b00000000000000000000111000101001;
			12'b11101010 		: log = 32'b00000000000000000000111000111000;
			12'b11101011 		: log = 32'b00000000000000000000111001001000;
			12'b11101100 		: log = 32'b00000000000000000000111001010111;
			12'b11101101 		: log = 32'b00000000000000000000111001100110;
			12'b11101110 		: log = 32'b00000000000000000000111001110101;
			12'b11101111 		: log = 32'b00000000000000000000111010000100;
			12'b11110000 		: log = 32'b00000000000000000000111010010011;
			12'b11110001 		: log = 32'b00000000000000000000111010100010;
			12'b11110010 		: log = 32'b00000000000000000000111010110001;
			12'b11110011 		: log = 32'b00000000000000000000111011000001;
			12'b11110100 		: log = 32'b00000000000000000000111011010000;
			12'b11110101 		: log = 32'b00000000000000000000111011011111;
			12'b11110110 		: log = 32'b00000000000000000000111011101110;
			12'b11110111 		: log = 32'b00000000000000000000111011111101;
			12'b11111000 		: log = 32'b00000000000000000000111100001100;
			12'b11111001 		: log = 32'b00000000000000000000111100011011;
			12'b11111010 		: log = 32'b00000000000000000000111100101010;
			12'b11111011 		: log = 32'b00000000000000000000111100111001;
			12'b11111100 		: log = 32'b00000000000000000000111101001000;
			12'b11111101 		: log = 32'b00000000000000000000111101010111;
			12'b11111110 		: log = 32'b00000000000000000000111101100110;
			12'b11111111 		: log = 32'b00000000000000000000111101110110;
			12'b100000000 		: log = 32'b00000000000000000000111110000101;
			12'b100000001 		: log = 32'b00000000000000000000111110010100;
			12'b100000010 		: log = 32'b00000000000000000000111110100011;
			12'b100000011 		: log = 32'b00000000000000000000111110110010;
			12'b100000100 		: log = 32'b00000000000000000000111111000001;
			12'b100000101 		: log = 32'b00000000000000000000111111010000;
			12'b100000110 		: log = 32'b00000000000000000000111111011111;
			12'b100000111 		: log = 32'b00000000000000000000111111101110;
			12'b100001000 		: log = 32'b00000000000000000000111111111101;
			12'b100001001 		: log = 32'b00000000000000000001000000001100;
			12'b100001010 		: log = 32'b00000000000000000001000000011011;
			12'b100001011 		: log = 32'b00000000000000000001000000101010;
			12'b100001100 		: log = 32'b00000000000000000001000000111001;
			12'b100001101 		: log = 32'b00000000000000000001000001001000;
			12'b100001110 		: log = 32'b00000000000000000001000001010111;
			12'b100001111 		: log = 32'b00000000000000000001000001100110;
			12'b100010000 		: log = 32'b00000000000000000001000001110101;
			12'b100010001 		: log = 32'b00000000000000000001000010000100;
			12'b100010010 		: log = 32'b00000000000000000001000010010011;
			12'b100010011 		: log = 32'b00000000000000000001000010100010;
			12'b100010100 		: log = 32'b00000000000000000001000010110001;
			12'b100010101 		: log = 32'b00000000000000000001000011000000;
			12'b100010110 		: log = 32'b00000000000000000001000011001111;
			12'b100010111 		: log = 32'b00000000000000000001000011011110;
			12'b100011000 		: log = 32'b00000000000000000001000011101101;
			12'b100011001 		: log = 32'b00000000000000000001000011111100;
			12'b100011010 		: log = 32'b00000000000000000001000100001011;
			12'b100011011 		: log = 32'b00000000000000000001000100011010;
			12'b100011100 		: log = 32'b00000000000000000001000100101001;
			12'b100011101 		: log = 32'b00000000000000000001000100111000;
			12'b100011110 		: log = 32'b00000000000000000001000101000111;
			12'b100011111 		: log = 32'b00000000000000000001000101010110;
			12'b100100000 		: log = 32'b00000000000000000001000101100101;
			12'b100100001 		: log = 32'b00000000000000000001000101110100;
			12'b100100010 		: log = 32'b00000000000000000001000110000011;
			12'b100100011 		: log = 32'b00000000000000000001000110010010;
			12'b100100100 		: log = 32'b00000000000000000001000110100000;
			12'b100100101 		: log = 32'b00000000000000000001000110101111;
			12'b100100110 		: log = 32'b00000000000000000001000110111110;
			12'b100100111 		: log = 32'b00000000000000000001000111001101;
			12'b100101000 		: log = 32'b00000000000000000001000111011100;
			12'b100101001 		: log = 32'b00000000000000000001000111101011;
			12'b100101010 		: log = 32'b00000000000000000001000111111010;
			12'b100101011 		: log = 32'b00000000000000000001001000001001;
			12'b100101100 		: log = 32'b00000000000000000001001000011000;
			12'b100101101 		: log = 32'b00000000000000000001001000100111;
			12'b100101110 		: log = 32'b00000000000000000001001000110110;
			12'b100101111 		: log = 32'b00000000000000000001001001000101;
			12'b100110000 		: log = 32'b00000000000000000001001001010011;
			12'b100110001 		: log = 32'b00000000000000000001001001100010;
			12'b100110010 		: log = 32'b00000000000000000001001001110001;
			12'b100110011 		: log = 32'b00000000000000000001001010000000;
			12'b100110100 		: log = 32'b00000000000000000001001010001111;
			12'b100110101 		: log = 32'b00000000000000000001001010011110;
			12'b100110110 		: log = 32'b00000000000000000001001010101101;
			12'b100110111 		: log = 32'b00000000000000000001001010111100;
			12'b100111000 		: log = 32'b00000000000000000001001011001011;
			12'b100111001 		: log = 32'b00000000000000000001001011011001;
			12'b100111010 		: log = 32'b00000000000000000001001011101000;
			12'b100111011 		: log = 32'b00000000000000000001001011110111;
			12'b100111100 		: log = 32'b00000000000000000001001100000110;
			12'b100111101 		: log = 32'b00000000000000000001001100010101;
			12'b100111110 		: log = 32'b00000000000000000001001100100100;
			12'b100111111 		: log = 32'b00000000000000000001001100110010;
			12'b101000000 		: log = 32'b00000000000000000001001101000001;
			12'b101000001 		: log = 32'b00000000000000000001001101010000;
			12'b101000010 		: log = 32'b00000000000000000001001101011111;
			12'b101000011 		: log = 32'b00000000000000000001001101101110;
			12'b101000100 		: log = 32'b00000000000000000001001101111101;
			12'b101000101 		: log = 32'b00000000000000000001001110001100;
			12'b101000110 		: log = 32'b00000000000000000001001110011010;
			12'b101000111 		: log = 32'b00000000000000000001001110101001;
			12'b101001000 		: log = 32'b00000000000000000001001110111000;
			12'b101001001 		: log = 32'b00000000000000000001001111000111;
			12'b101001010 		: log = 32'b00000000000000000001001111010110;
			12'b101001011 		: log = 32'b00000000000000000001001111100100;
			12'b101001100 		: log = 32'b00000000000000000001001111110011;
			12'b101001101 		: log = 32'b00000000000000000001010000000010;
			12'b101001110 		: log = 32'b00000000000000000001010000010001;
			12'b101001111 		: log = 32'b00000000000000000001010000100000;
			12'b101010000 		: log = 32'b00000000000000000001010000101110;
			12'b101010001 		: log = 32'b00000000000000000001010000111101;
			12'b101010010 		: log = 32'b00000000000000000001010001001100;
			12'b101010011 		: log = 32'b00000000000000000001010001011011;
			12'b101010100 		: log = 32'b00000000000000000001010001101001;
			12'b101010101 		: log = 32'b00000000000000000001010001111000;
			12'b101010110 		: log = 32'b00000000000000000001010010000111;
			12'b101010111 		: log = 32'b00000000000000000001010010010110;
			12'b101011000 		: log = 32'b00000000000000000001010010100101;
			12'b101011001 		: log = 32'b00000000000000000001010010110011;
			12'b101011010 		: log = 32'b00000000000000000001010011000010;
			12'b101011011 		: log = 32'b00000000000000000001010011010001;
			12'b101011100 		: log = 32'b00000000000000000001010011100000;
			12'b101011101 		: log = 32'b00000000000000000001010011101110;
			12'b101011110 		: log = 32'b00000000000000000001010011111101;
			12'b101011111 		: log = 32'b00000000000000000001010100001100;
			12'b101100000 		: log = 32'b00000000000000000001010100011011;
			12'b101100001 		: log = 32'b00000000000000000001010100101001;
			12'b101100010 		: log = 32'b00000000000000000001010100111000;
			12'b101100011 		: log = 32'b00000000000000000001010101000111;
			12'b101100100 		: log = 32'b00000000000000000001010101010101;
			12'b101100101 		: log = 32'b00000000000000000001010101100100;
			12'b101100110 		: log = 32'b00000000000000000001010101110011;
			12'b101100111 		: log = 32'b00000000000000000001010110000010;
			12'b101101000 		: log = 32'b00000000000000000001010110010000;
			12'b101101001 		: log = 32'b00000000000000000001010110011111;
			12'b101101010 		: log = 32'b00000000000000000001010110101110;
			12'b101101011 		: log = 32'b00000000000000000001010110111100;
			12'b101101100 		: log = 32'b00000000000000000001010111001011;
			12'b101101101 		: log = 32'b00000000000000000001010111011010;
			12'b101101110 		: log = 32'b00000000000000000001010111101000;
			12'b101101111 		: log = 32'b00000000000000000001010111110111;
			12'b101110000 		: log = 32'b00000000000000000001011000000110;
			12'b101110001 		: log = 32'b00000000000000000001011000010101;
			12'b101110010 		: log = 32'b00000000000000000001011000100011;
			12'b101110011 		: log = 32'b00000000000000000001011000110010;
			12'b101110100 		: log = 32'b00000000000000000001011001000001;
			12'b101110101 		: log = 32'b00000000000000000001011001001111;
			12'b101110110 		: log = 32'b00000000000000000001011001011110;
			12'b101110111 		: log = 32'b00000000000000000001011001101101;
			12'b101111000 		: log = 32'b00000000000000000001011001111011;
			12'b101111001 		: log = 32'b00000000000000000001011010001010;
			12'b101111010 		: log = 32'b00000000000000000001011010011000;
			12'b101111011 		: log = 32'b00000000000000000001011010100111;
			12'b101111100 		: log = 32'b00000000000000000001011010110110;
			12'b101111101 		: log = 32'b00000000000000000001011011000100;
			12'b101111110 		: log = 32'b00000000000000000001011011010011;
			12'b101111111 		: log = 32'b00000000000000000001011011100010;
			12'b110000000 		: log = 32'b00000000000000000001011011110000;
			12'b110000001 		: log = 32'b00000000000000000001011011111111;
			12'b110000010 		: log = 32'b00000000000000000001011100001110;
			12'b110000011 		: log = 32'b00000000000000000001011100011100;
			12'b110000100 		: log = 32'b00000000000000000001011100101011;
			12'b110000101 		: log = 32'b00000000000000000001011100111001;
			12'b110000110 		: log = 32'b00000000000000000001011101001000;
			12'b110000111 		: log = 32'b00000000000000000001011101010111;
			12'b110001000 		: log = 32'b00000000000000000001011101100101;
			12'b110001001 		: log = 32'b00000000000000000001011101110100;
			12'b110001010 		: log = 32'b00000000000000000001011110000010;
			12'b110001011 		: log = 32'b00000000000000000001011110010001;
			12'b110001100 		: log = 32'b00000000000000000001011110100000;
			12'b110001101 		: log = 32'b00000000000000000001011110101110;
			12'b110001110 		: log = 32'b00000000000000000001011110111101;
			12'b110001111 		: log = 32'b00000000000000000001011111001011;
			12'b110010000 		: log = 32'b00000000000000000001011111011010;
			12'b110010001 		: log = 32'b00000000000000000001011111101001;
			12'b110010010 		: log = 32'b00000000000000000001011111110111;
			12'b110010011 		: log = 32'b00000000000000000001100000000110;
			12'b110010100 		: log = 32'b00000000000000000001100000010100;
			12'b110010101 		: log = 32'b00000000000000000001100000100011;
			12'b110010110 		: log = 32'b00000000000000000001100000110001;
			12'b110010111 		: log = 32'b00000000000000000001100001000000;
			12'b110011000 		: log = 32'b00000000000000000001100001001110;
			12'b110011001 		: log = 32'b00000000000000000001100001011101;
			12'b110011010 		: log = 32'b00000000000000000001100001101100;
			12'b110011011 		: log = 32'b00000000000000000001100001111010;
			12'b110011100 		: log = 32'b00000000000000000001100010001001;
			12'b110011101 		: log = 32'b00000000000000000001100010010111;
			12'b110011110 		: log = 32'b00000000000000000001100010100110;
			12'b110011111 		: log = 32'b00000000000000000001100010110100;
			12'b110100000 		: log = 32'b00000000000000000001100011000011;
			12'b110100001 		: log = 32'b00000000000000000001100011010001;
			12'b110100010 		: log = 32'b00000000000000000001100011100000;
			12'b110100011 		: log = 32'b00000000000000000001100011101110;
			12'b110100100 		: log = 32'b00000000000000000001100011111101;
			12'b110100101 		: log = 32'b00000000000000000001100100001011;
			12'b110100110 		: log = 32'b00000000000000000001100100011010;
			12'b110100111 		: log = 32'b00000000000000000001100100101000;
			12'b110101000 		: log = 32'b00000000000000000001100100110111;
			12'b110101001 		: log = 32'b00000000000000000001100101000101;
			12'b110101010 		: log = 32'b00000000000000000001100101010100;
			12'b110101011 		: log = 32'b00000000000000000001100101100010;
			12'b110101100 		: log = 32'b00000000000000000001100101110001;
			12'b110101101 		: log = 32'b00000000000000000001100101111111;
			12'b110101110 		: log = 32'b00000000000000000001100110001110;
			12'b110101111 		: log = 32'b00000000000000000001100110011100;
			12'b110110000 		: log = 32'b00000000000000000001100110101011;
			12'b110110001 		: log = 32'b00000000000000000001100110111001;
			12'b110110010 		: log = 32'b00000000000000000001100111001000;
			12'b110110011 		: log = 32'b00000000000000000001100111010110;
			12'b110110100 		: log = 32'b00000000000000000001100111100101;
			12'b110110101 		: log = 32'b00000000000000000001100111110011;
			12'b110110110 		: log = 32'b00000000000000000001101000000010;
			12'b110110111 		: log = 32'b00000000000000000001101000010000;
			12'b110111000 		: log = 32'b00000000000000000001101000011110;
			12'b110111001 		: log = 32'b00000000000000000001101000101101;
			12'b110111010 		: log = 32'b00000000000000000001101000111011;
			12'b110111011 		: log = 32'b00000000000000000001101001001010;
			12'b110111100 		: log = 32'b00000000000000000001101001011000;
			12'b110111101 		: log = 32'b00000000000000000001101001100111;
			12'b110111110 		: log = 32'b00000000000000000001101001110101;
			12'b110111111 		: log = 32'b00000000000000000001101010000100;
			12'b111000000 		: log = 32'b00000000000000000001101010010010;
			12'b111000001 		: log = 32'b00000000000000000001101010100000;
			12'b111000010 		: log = 32'b00000000000000000001101010101111;
			12'b111000011 		: log = 32'b00000000000000000001101010111101;
			12'b111000100 		: log = 32'b00000000000000000001101011001100;
			12'b111000101 		: log = 32'b00000000000000000001101011011010;
			12'b111000110 		: log = 32'b00000000000000000001101011101000;
			12'b111000111 		: log = 32'b00000000000000000001101011110111;
			12'b111001000 		: log = 32'b00000000000000000001101100000101;
			12'b111001001 		: log = 32'b00000000000000000001101100010100;
			12'b111001010 		: log = 32'b00000000000000000001101100100010;
			12'b111001011 		: log = 32'b00000000000000000001101100110000;
			12'b111001100 		: log = 32'b00000000000000000001101100111111;
			12'b111001101 		: log = 32'b00000000000000000001101101001101;
			12'b111001110 		: log = 32'b00000000000000000001101101011100;
			12'b111001111 		: log = 32'b00000000000000000001101101101010;
			12'b111010000 		: log = 32'b00000000000000000001101101111000;
			12'b111010001 		: log = 32'b00000000000000000001101110000111;
			12'b111010010 		: log = 32'b00000000000000000001101110010101;
			12'b111010011 		: log = 32'b00000000000000000001101110100011;
			12'b111010100 		: log = 32'b00000000000000000001101110110010;
			12'b111010101 		: log = 32'b00000000000000000001101111000000;
			12'b111010110 		: log = 32'b00000000000000000001101111001110;
			12'b111010111 		: log = 32'b00000000000000000001101111011101;
			12'b111011000 		: log = 32'b00000000000000000001101111101011;
			12'b111011001 		: log = 32'b00000000000000000001101111111010;
			12'b111011010 		: log = 32'b00000000000000000001110000001000;
			12'b111011011 		: log = 32'b00000000000000000001110000010110;
			12'b111011100 		: log = 32'b00000000000000000001110000100101;
			12'b111011101 		: log = 32'b00000000000000000001110000110011;
			12'b111011110 		: log = 32'b00000000000000000001110001000001;
			12'b111011111 		: log = 32'b00000000000000000001110001010000;
			12'b111100000 		: log = 32'b00000000000000000001110001011110;
			12'b111100001 		: log = 32'b00000000000000000001110001101100;
			12'b111100010 		: log = 32'b00000000000000000001110001111010;
			12'b111100011 		: log = 32'b00000000000000000001110010001001;
			12'b111100100 		: log = 32'b00000000000000000001110010010111;
			12'b111100101 		: log = 32'b00000000000000000001110010100101;
			12'b111100110 		: log = 32'b00000000000000000001110010110100;
			12'b111100111 		: log = 32'b00000000000000000001110011000010;
			12'b111101000 		: log = 32'b00000000000000000001110011010000;
			12'b111101001 		: log = 32'b00000000000000000001110011011111;
			12'b111101010 		: log = 32'b00000000000000000001110011101101;
			12'b111101011 		: log = 32'b00000000000000000001110011111011;
			12'b111101100 		: log = 32'b00000000000000000001110100001001;
			12'b111101101 		: log = 32'b00000000000000000001110100011000;
			12'b111101110 		: log = 32'b00000000000000000001110100100110;
			12'b111101111 		: log = 32'b00000000000000000001110100110100;
			12'b111110000 		: log = 32'b00000000000000000001110101000011;
			12'b111110001 		: log = 32'b00000000000000000001110101010001;
			12'b111110010 		: log = 32'b00000000000000000001110101011111;
			12'b111110011 		: log = 32'b00000000000000000001110101101101;
			12'b111110100 		: log = 32'b00000000000000000001110101111100;
			12'b111110101 		: log = 32'b00000000000000000001110110001010;
			12'b111110110 		: log = 32'b00000000000000000001110110011000;
			12'b111110111 		: log = 32'b00000000000000000001110110100110;
			12'b111111000 		: log = 32'b00000000000000000001110110110101;
			12'b111111001 		: log = 32'b00000000000000000001110111000011;
			12'b111111010 		: log = 32'b00000000000000000001110111010001;
			12'b111111011 		: log = 32'b00000000000000000001110111011111;
			12'b111111100 		: log = 32'b00000000000000000001110111101110;
			12'b111111101 		: log = 32'b00000000000000000001110111111100;
			12'b111111110 		: log = 32'b00000000000000000001111000001010;
			12'b111111111 		: log = 32'b00000000000000000001111000011000;
			12'b1000000000 		: log = 32'b00000000000000000001111000100111;
			12'b1000000001 		: log = 32'b00000000000000000001111000110101;
			12'b1000000010 		: log = 32'b00000000000000000001111001000011;
			12'b1000000011 		: log = 32'b00000000000000000001111001010001;
			12'b1000000100 		: log = 32'b00000000000000000001111001011111;
			12'b1000000101 		: log = 32'b00000000000000000001111001101110;
			12'b1000000110 		: log = 32'b00000000000000000001111001111100;
			12'b1000000111 		: log = 32'b00000000000000000001111010001010;
			12'b1000001000 		: log = 32'b00000000000000000001111010011000;
			12'b1000001001 		: log = 32'b00000000000000000001111010100110;
			12'b1000001010 		: log = 32'b00000000000000000001111010110101;
			12'b1000001011 		: log = 32'b00000000000000000001111011000011;
			12'b1000001100 		: log = 32'b00000000000000000001111011010001;
			12'b1000001101 		: log = 32'b00000000000000000001111011011111;
			12'b1000001110 		: log = 32'b00000000000000000001111011101101;
			12'b1000001111 		: log = 32'b00000000000000000001111011111100;
			12'b1000010000 		: log = 32'b00000000000000000001111100001010;
			12'b1000010001 		: log = 32'b00000000000000000001111100011000;
			12'b1000010010 		: log = 32'b00000000000000000001111100100110;
			12'b1000010011 		: log = 32'b00000000000000000001111100110100;
			12'b1000010100 		: log = 32'b00000000000000000001111101000010;
			12'b1000010101 		: log = 32'b00000000000000000001111101010001;
			12'b1000010110 		: log = 32'b00000000000000000001111101011111;
			12'b1000010111 		: log = 32'b00000000000000000001111101101101;
			12'b1000011000 		: log = 32'b00000000000000000001111101111011;
			12'b1000011001 		: log = 32'b00000000000000000001111110001001;
			12'b1000011010 		: log = 32'b00000000000000000001111110010111;
			12'b1000011011 		: log = 32'b00000000000000000001111110100101;
			12'b1000011100 		: log = 32'b00000000000000000001111110110100;
			12'b1000011101 		: log = 32'b00000000000000000001111111000010;
			12'b1000011110 		: log = 32'b00000000000000000001111111010000;
			12'b1000011111 		: log = 32'b00000000000000000001111111011110;
			12'b1000100000 		: log = 32'b00000000000000000001111111101100;
			12'b1000100001 		: log = 32'b00000000000000000001111111111010;
			12'b1000100010 		: log = 32'b00000000000000000010000000001000;
			12'b1000100011 		: log = 32'b00000000000000000010000000010110;
			12'b1000100100 		: log = 32'b00000000000000000010000000100101;
			12'b1000100101 		: log = 32'b00000000000000000010000000110011;
			12'b1000100110 		: log = 32'b00000000000000000010000001000001;
			12'b1000100111 		: log = 32'b00000000000000000010000001001111;
			12'b1000101000 		: log = 32'b00000000000000000010000001011101;
			12'b1000101001 		: log = 32'b00000000000000000010000001101011;
			12'b1000101010 		: log = 32'b00000000000000000010000001111001;
			12'b1000101011 		: log = 32'b00000000000000000010000010000111;
			12'b1000101100 		: log = 32'b00000000000000000010000010010101;
			12'b1000101101 		: log = 32'b00000000000000000010000010100011;
			12'b1000101110 		: log = 32'b00000000000000000010000010110010;
			12'b1000101111 		: log = 32'b00000000000000000010000011000000;
			12'b1000110000 		: log = 32'b00000000000000000010000011001110;
			12'b1000110001 		: log = 32'b00000000000000000010000011011100;
			12'b1000110010 		: log = 32'b00000000000000000010000011101010;
			12'b1000110011 		: log = 32'b00000000000000000010000011111000;
			12'b1000110100 		: log = 32'b00000000000000000010000100000110;
			12'b1000110101 		: log = 32'b00000000000000000010000100010100;
			12'b1000110110 		: log = 32'b00000000000000000010000100100010;
			12'b1000110111 		: log = 32'b00000000000000000010000100110000;
			12'b1000111000 		: log = 32'b00000000000000000010000100111110;
			12'b1000111001 		: log = 32'b00000000000000000010000101001100;
			12'b1000111010 		: log = 32'b00000000000000000010000101011010;
			12'b1000111011 		: log = 32'b00000000000000000010000101101000;
			12'b1000111100 		: log = 32'b00000000000000000010000101110110;
			12'b1000111101 		: log = 32'b00000000000000000010000110000100;
			12'b1000111110 		: log = 32'b00000000000000000010000110010010;
			12'b1000111111 		: log = 32'b00000000000000000010000110100000;
			12'b1001000000 		: log = 32'b00000000000000000010000110101110;
			12'b1001000001 		: log = 32'b00000000000000000010000110111101;
			12'b1001000010 		: log = 32'b00000000000000000010000111001011;
			12'b1001000011 		: log = 32'b00000000000000000010000111011001;
			12'b1001000100 		: log = 32'b00000000000000000010000111100111;
			12'b1001000101 		: log = 32'b00000000000000000010000111110101;
			12'b1001000110 		: log = 32'b00000000000000000010001000000011;
			12'b1001000111 		: log = 32'b00000000000000000010001000010001;
			12'b1001001000 		: log = 32'b00000000000000000010001000011111;
			12'b1001001001 		: log = 32'b00000000000000000010001000101101;
			12'b1001001010 		: log = 32'b00000000000000000010001000111011;
			12'b1001001011 		: log = 32'b00000000000000000010001001001001;
			12'b1001001100 		: log = 32'b00000000000000000010001001010111;
			12'b1001001101 		: log = 32'b00000000000000000010001001100101;
			12'b1001001110 		: log = 32'b00000000000000000010001001110011;
			12'b1001001111 		: log = 32'b00000000000000000010001010000001;
			12'b1001010000 		: log = 32'b00000000000000000010001010001111;
			12'b1001010001 		: log = 32'b00000000000000000010001010011101;
			12'b1001010010 		: log = 32'b00000000000000000010001010101010;
			12'b1001010011 		: log = 32'b00000000000000000010001010111000;
			12'b1001010100 		: log = 32'b00000000000000000010001011000110;
			12'b1001010101 		: log = 32'b00000000000000000010001011010100;
			12'b1001010110 		: log = 32'b00000000000000000010001011100010;
			12'b1001010111 		: log = 32'b00000000000000000010001011110000;
			12'b1001011000 		: log = 32'b00000000000000000010001011111110;
			12'b1001011001 		: log = 32'b00000000000000000010001100001100;
			12'b1001011010 		: log = 32'b00000000000000000010001100011010;
			12'b1001011011 		: log = 32'b00000000000000000010001100101000;
			12'b1001011100 		: log = 32'b00000000000000000010001100110110;
			12'b1001011101 		: log = 32'b00000000000000000010001101000100;
			12'b1001011110 		: log = 32'b00000000000000000010001101010010;
			12'b1001011111 		: log = 32'b00000000000000000010001101100000;
			12'b1001100000 		: log = 32'b00000000000000000010001101101110;
			12'b1001100001 		: log = 32'b00000000000000000010001101111100;
			12'b1001100010 		: log = 32'b00000000000000000010001110001010;
			12'b1001100011 		: log = 32'b00000000000000000010001110011000;
			12'b1001100100 		: log = 32'b00000000000000000010001110100110;
			12'b1001100101 		: log = 32'b00000000000000000010001110110011;
			12'b1001100110 		: log = 32'b00000000000000000010001111000001;
			12'b1001100111 		: log = 32'b00000000000000000010001111001111;
			12'b1001101000 		: log = 32'b00000000000000000010001111011101;
			12'b1001101001 		: log = 32'b00000000000000000010001111101011;
			12'b1001101010 		: log = 32'b00000000000000000010001111111001;
			12'b1001101011 		: log = 32'b00000000000000000010010000000111;
			12'b1001101100 		: log = 32'b00000000000000000010010000010101;
			12'b1001101101 		: log = 32'b00000000000000000010010000100011;
			12'b1001101110 		: log = 32'b00000000000000000010010000110001;
			12'b1001101111 		: log = 32'b00000000000000000010010000111110;
			12'b1001110000 		: log = 32'b00000000000000000010010001001100;
			12'b1001110001 		: log = 32'b00000000000000000010010001011010;
			12'b1001110010 		: log = 32'b00000000000000000010010001101000;
			12'b1001110011 		: log = 32'b00000000000000000010010001110110;
			12'b1001110100 		: log = 32'b00000000000000000010010010000100;
			12'b1001110101 		: log = 32'b00000000000000000010010010010010;
			12'b1001110110 		: log = 32'b00000000000000000010010010100000;
			12'b1001110111 		: log = 32'b00000000000000000010010010101101;
			12'b1001111000 		: log = 32'b00000000000000000010010010111011;
			12'b1001111001 		: log = 32'b00000000000000000010010011001001;
			12'b1001111010 		: log = 32'b00000000000000000010010011010111;
			12'b1001111011 		: log = 32'b00000000000000000010010011100101;
			12'b1001111100 		: log = 32'b00000000000000000010010011110011;
			12'b1001111101 		: log = 32'b00000000000000000010010100000001;
			12'b1001111110 		: log = 32'b00000000000000000010010100001110;
			12'b1001111111 		: log = 32'b00000000000000000010010100011100;
			12'b1010000000 		: log = 32'b00000000000000000010010100101010;
			12'b1010000001 		: log = 32'b00000000000000000010010100111000;
			12'b1010000010 		: log = 32'b00000000000000000010010101000110;
			12'b1010000011 		: log = 32'b00000000000000000010010101010100;
			12'b1010000100 		: log = 32'b00000000000000000010010101100001;
			12'b1010000101 		: log = 32'b00000000000000000010010101101111;
			12'b1010000110 		: log = 32'b00000000000000000010010101111101;
			12'b1010000111 		: log = 32'b00000000000000000010010110001011;
			12'b1010001000 		: log = 32'b00000000000000000010010110011001;
			12'b1010001001 		: log = 32'b00000000000000000010010110100111;
			12'b1010001010 		: log = 32'b00000000000000000010010110110100;
			12'b1010001011 		: log = 32'b00000000000000000010010111000010;
			12'b1010001100 		: log = 32'b00000000000000000010010111010000;
			12'b1010001101 		: log = 32'b00000000000000000010010111011110;
			12'b1010001110 		: log = 32'b00000000000000000010010111101100;
			12'b1010001111 		: log = 32'b00000000000000000010010111111001;
			12'b1010010000 		: log = 32'b00000000000000000010011000000111;
			12'b1010010001 		: log = 32'b00000000000000000010011000010101;
			12'b1010010010 		: log = 32'b00000000000000000010011000100011;
			12'b1010010011 		: log = 32'b00000000000000000010011000110001;
			12'b1010010100 		: log = 32'b00000000000000000010011000111110;
			12'b1010010101 		: log = 32'b00000000000000000010011001001100;
			12'b1010010110 		: log = 32'b00000000000000000010011001011010;
			12'b1010010111 		: log = 32'b00000000000000000010011001101000;
			12'b1010011000 		: log = 32'b00000000000000000010011001110101;
			12'b1010011001 		: log = 32'b00000000000000000010011010000011;
			12'b1010011010 		: log = 32'b00000000000000000010011010010001;
			12'b1010011011 		: log = 32'b00000000000000000010011010011111;
			12'b1010011100 		: log = 32'b00000000000000000010011010101100;
			12'b1010011101 		: log = 32'b00000000000000000010011010111010;
			12'b1010011110 		: log = 32'b00000000000000000010011011001000;
			12'b1010011111 		: log = 32'b00000000000000000010011011010110;
			12'b1010100000 		: log = 32'b00000000000000000010011011100011;
			12'b1010100001 		: log = 32'b00000000000000000010011011110001;
			12'b1010100010 		: log = 32'b00000000000000000010011011111111;
			12'b1010100011 		: log = 32'b00000000000000000010011100001101;
			12'b1010100100 		: log = 32'b00000000000000000010011100011010;
			12'b1010100101 		: log = 32'b00000000000000000010011100101000;
			12'b1010100110 		: log = 32'b00000000000000000010011100110110;
			12'b1010100111 		: log = 32'b00000000000000000010011101000100;
			12'b1010101000 		: log = 32'b00000000000000000010011101010001;
			12'b1010101001 		: log = 32'b00000000000000000010011101011111;
			12'b1010101010 		: log = 32'b00000000000000000010011101101101;
			12'b1010101011 		: log = 32'b00000000000000000010011101111010;
			12'b1010101100 		: log = 32'b00000000000000000010011110001000;
			12'b1010101101 		: log = 32'b00000000000000000010011110010110;
			12'b1010101110 		: log = 32'b00000000000000000010011110100100;
			12'b1010101111 		: log = 32'b00000000000000000010011110110001;
			12'b1010110000 		: log = 32'b00000000000000000010011110111111;
			12'b1010110001 		: log = 32'b00000000000000000010011111001101;
			12'b1010110010 		: log = 32'b00000000000000000010011111011010;
			12'b1010110011 		: log = 32'b00000000000000000010011111101000;
			12'b1010110100 		: log = 32'b00000000000000000010011111110110;
			12'b1010110101 		: log = 32'b00000000000000000010100000000011;
			12'b1010110110 		: log = 32'b00000000000000000010100000010001;
			12'b1010110111 		: log = 32'b00000000000000000010100000011111;
			12'b1010111000 		: log = 32'b00000000000000000010100000101101;
			12'b1010111001 		: log = 32'b00000000000000000010100000111010;
			12'b1010111010 		: log = 32'b00000000000000000010100001001000;
			12'b1010111011 		: log = 32'b00000000000000000010100001010110;
			12'b1010111100 		: log = 32'b00000000000000000010100001100011;
			12'b1010111101 		: log = 32'b00000000000000000010100001110001;
			12'b1010111110 		: log = 32'b00000000000000000010100001111111;
			12'b1010111111 		: log = 32'b00000000000000000010100010001100;
			12'b1011000000 		: log = 32'b00000000000000000010100010011010;
			12'b1011000001 		: log = 32'b00000000000000000010100010100111;
			12'b1011000010 		: log = 32'b00000000000000000010100010110101;
			12'b1011000011 		: log = 32'b00000000000000000010100011000011;
			12'b1011000100 		: log = 32'b00000000000000000010100011010000;
			12'b1011000101 		: log = 32'b00000000000000000010100011011110;
			12'b1011000110 		: log = 32'b00000000000000000010100011101100;
			12'b1011000111 		: log = 32'b00000000000000000010100011111001;
			12'b1011001000 		: log = 32'b00000000000000000010100100000111;
			12'b1011001001 		: log = 32'b00000000000000000010100100010101;
			12'b1011001010 		: log = 32'b00000000000000000010100100100010;
			12'b1011001011 		: log = 32'b00000000000000000010100100110000;
			12'b1011001100 		: log = 32'b00000000000000000010100100111101;
			12'b1011001101 		: log = 32'b00000000000000000010100101001011;
			12'b1011001110 		: log = 32'b00000000000000000010100101011001;
			12'b1011001111 		: log = 32'b00000000000000000010100101100110;
			12'b1011010000 		: log = 32'b00000000000000000010100101110100;
			12'b1011010001 		: log = 32'b00000000000000000010100110000010;
			12'b1011010010 		: log = 32'b00000000000000000010100110001111;
			12'b1011010011 		: log = 32'b00000000000000000010100110011101;
			12'b1011010100 		: log = 32'b00000000000000000010100110101010;
			12'b1011010101 		: log = 32'b00000000000000000010100110111000;
			12'b1011010110 		: log = 32'b00000000000000000010100111000110;
			12'b1011010111 		: log = 32'b00000000000000000010100111010011;
			12'b1011011000 		: log = 32'b00000000000000000010100111100001;
			12'b1011011001 		: log = 32'b00000000000000000010100111101110;
			12'b1011011010 		: log = 32'b00000000000000000010100111111100;
			12'b1011011011 		: log = 32'b00000000000000000010101000001001;
			12'b1011011100 		: log = 32'b00000000000000000010101000010111;
			12'b1011011101 		: log = 32'b00000000000000000010101000100101;
			12'b1011011110 		: log = 32'b00000000000000000010101000110010;
			12'b1011011111 		: log = 32'b00000000000000000010101001000000;
			12'b1011100000 		: log = 32'b00000000000000000010101001001101;
			12'b1011100001 		: log = 32'b00000000000000000010101001011011;
			12'b1011100010 		: log = 32'b00000000000000000010101001101000;
			12'b1011100011 		: log = 32'b00000000000000000010101001110110;
			12'b1011100100 		: log = 32'b00000000000000000010101010000100;
			12'b1011100101 		: log = 32'b00000000000000000010101010010001;
			12'b1011100110 		: log = 32'b00000000000000000010101010011111;
			12'b1011100111 		: log = 32'b00000000000000000010101010101100;
			12'b1011101000 		: log = 32'b00000000000000000010101010111010;
			12'b1011101001 		: log = 32'b00000000000000000010101011000111;
			12'b1011101010 		: log = 32'b00000000000000000010101011010101;
			12'b1011101011 		: log = 32'b00000000000000000010101011100010;
			12'b1011101100 		: log = 32'b00000000000000000010101011110000;
			12'b1011101101 		: log = 32'b00000000000000000010101011111101;
			12'b1011101110 		: log = 32'b00000000000000000010101100001011;
			12'b1011101111 		: log = 32'b00000000000000000010101100011000;
			12'b1011110000 		: log = 32'b00000000000000000010101100100110;
			12'b1011110001 		: log = 32'b00000000000000000010101100110011;
			12'b1011110010 		: log = 32'b00000000000000000010101101000001;
			12'b1011110011 		: log = 32'b00000000000000000010101101001110;
			12'b1011110100 		: log = 32'b00000000000000000010101101011100;
			12'b1011110101 		: log = 32'b00000000000000000010101101101010;
			12'b1011110110 		: log = 32'b00000000000000000010101101110111;
			12'b1011110111 		: log = 32'b00000000000000000010101110000101;
			12'b1011111000 		: log = 32'b00000000000000000010101110010010;
			12'b1011111001 		: log = 32'b00000000000000000010101110011111;
			12'b1011111010 		: log = 32'b00000000000000000010101110101101;
			12'b1011111011 		: log = 32'b00000000000000000010101110111010;
			12'b1011111100 		: log = 32'b00000000000000000010101111001000;
			12'b1011111101 		: log = 32'b00000000000000000010101111010101;
			12'b1011111110 		: log = 32'b00000000000000000010101111100011;
			12'b1011111111 		: log = 32'b00000000000000000010101111110000;
			12'b1100000000 		: log = 32'b00000000000000000010101111111110;
			12'b1100000001 		: log = 32'b00000000000000000010110000001011;
			12'b1100000010 		: log = 32'b00000000000000000010110000011001;
			12'b1100000011 		: log = 32'b00000000000000000010110000100110;
			12'b1100000100 		: log = 32'b00000000000000000010110000110100;
			12'b1100000101 		: log = 32'b00000000000000000010110001000001;
			12'b1100000110 		: log = 32'b00000000000000000010110001001111;
			12'b1100000111 		: log = 32'b00000000000000000010110001011100;
			12'b1100001000 		: log = 32'b00000000000000000010110001101010;
			12'b1100001001 		: log = 32'b00000000000000000010110001110111;
			12'b1100001010 		: log = 32'b00000000000000000010110010000100;
			12'b1100001011 		: log = 32'b00000000000000000010110010010010;
			12'b1100001100 		: log = 32'b00000000000000000010110010011111;
			12'b1100001101 		: log = 32'b00000000000000000010110010101101;
			12'b1100001110 		: log = 32'b00000000000000000010110010111010;
			12'b1100001111 		: log = 32'b00000000000000000010110011001000;
			12'b1100010000 		: log = 32'b00000000000000000010110011010101;
			12'b1100010001 		: log = 32'b00000000000000000010110011100011;
			12'b1100010010 		: log = 32'b00000000000000000010110011110000;
			12'b1100010011 		: log = 32'b00000000000000000010110011111101;
			12'b1100010100 		: log = 32'b00000000000000000010110100001011;
			12'b1100010101 		: log = 32'b00000000000000000010110100011000;
			12'b1100010110 		: log = 32'b00000000000000000010110100100110;
			12'b1100010111 		: log = 32'b00000000000000000010110100110011;
			12'b1100011000 		: log = 32'b00000000000000000010110101000000;
			12'b1100011001 		: log = 32'b00000000000000000010110101001110;
			12'b1100011010 		: log = 32'b00000000000000000010110101011011;
			12'b1100011011 		: log = 32'b00000000000000000010110101101001;
			12'b1100011100 		: log = 32'b00000000000000000010110101110110;
			12'b1100011101 		: log = 32'b00000000000000000010110110000011;
			12'b1100011110 		: log = 32'b00000000000000000010110110010001;
			12'b1100011111 		: log = 32'b00000000000000000010110110011110;
			12'b1100100000 		: log = 32'b00000000000000000010110110101100;
			12'b1100100001 		: log = 32'b00000000000000000010110110111001;
			12'b1100100010 		: log = 32'b00000000000000000010110111000110;
			12'b1100100011 		: log = 32'b00000000000000000010110111010100;
			12'b1100100100 		: log = 32'b00000000000000000010110111100001;
			12'b1100100101 		: log = 32'b00000000000000000010110111101111;
			12'b1100100110 		: log = 32'b00000000000000000010110111111100;
			12'b1100100111 		: log = 32'b00000000000000000010111000001001;
			12'b1100101000 		: log = 32'b00000000000000000010111000010111;
			12'b1100101001 		: log = 32'b00000000000000000010111000100100;
			12'b1100101010 		: log = 32'b00000000000000000010111000110001;
			12'b1100101011 		: log = 32'b00000000000000000010111000111111;
			12'b1100101100 		: log = 32'b00000000000000000010111001001100;
			12'b1100101101 		: log = 32'b00000000000000000010111001011001;
			12'b1100101110 		: log = 32'b00000000000000000010111001100111;
			12'b1100101111 		: log = 32'b00000000000000000010111001110100;
			12'b1100110000 		: log = 32'b00000000000000000010111010000001;
			12'b1100110001 		: log = 32'b00000000000000000010111010001111;
			12'b1100110010 		: log = 32'b00000000000000000010111010011100;
			12'b1100110011 		: log = 32'b00000000000000000010111010101001;
			12'b1100110100 		: log = 32'b00000000000000000010111010110111;
			12'b1100110101 		: log = 32'b00000000000000000010111011000100;
			12'b1100110110 		: log = 32'b00000000000000000010111011010001;
			12'b1100110111 		: log = 32'b00000000000000000010111011011111;
			12'b1100111000 		: log = 32'b00000000000000000010111011101100;
			12'b1100111001 		: log = 32'b00000000000000000010111011111001;
			12'b1100111010 		: log = 32'b00000000000000000010111100000111;
			12'b1100111011 		: log = 32'b00000000000000000010111100010100;
			12'b1100111100 		: log = 32'b00000000000000000010111100100001;
			12'b1100111101 		: log = 32'b00000000000000000010111100101111;
			12'b1100111110 		: log = 32'b00000000000000000010111100111100;
			12'b1100111111 		: log = 32'b00000000000000000010111101001001;
			12'b1101000000 		: log = 32'b00000000000000000010111101010111;
			12'b1101000001 		: log = 32'b00000000000000000010111101100100;
			12'b1101000010 		: log = 32'b00000000000000000010111101110001;
			12'b1101000011 		: log = 32'b00000000000000000010111101111110;
			12'b1101000100 		: log = 32'b00000000000000000010111110001100;
			12'b1101000101 		: log = 32'b00000000000000000010111110011001;
			12'b1101000110 		: log = 32'b00000000000000000010111110100110;
			12'b1101000111 		: log = 32'b00000000000000000010111110110100;
			12'b1101001000 		: log = 32'b00000000000000000010111111000001;
			12'b1101001001 		: log = 32'b00000000000000000010111111001110;
			12'b1101001010 		: log = 32'b00000000000000000010111111011011;
			12'b1101001011 		: log = 32'b00000000000000000010111111101001;
			12'b1101001100 		: log = 32'b00000000000000000010111111110110;
			12'b1101001101 		: log = 32'b00000000000000000011000000000011;
			12'b1101001110 		: log = 32'b00000000000000000011000000010000;
			12'b1101001111 		: log = 32'b00000000000000000011000000011110;
			12'b1101010000 		: log = 32'b00000000000000000011000000101011;
			12'b1101010001 		: log = 32'b00000000000000000011000000111000;
			12'b1101010010 		: log = 32'b00000000000000000011000001000110;
			12'b1101010011 		: log = 32'b00000000000000000011000001010011;
			12'b1101010100 		: log = 32'b00000000000000000011000001100000;
			12'b1101010101 		: log = 32'b00000000000000000011000001101101;
			12'b1101010110 		: log = 32'b00000000000000000011000001111010;
			12'b1101010111 		: log = 32'b00000000000000000011000010001000;
			12'b1101011000 		: log = 32'b00000000000000000011000010010101;
			12'b1101011001 		: log = 32'b00000000000000000011000010100010;
			12'b1101011010 		: log = 32'b00000000000000000011000010101111;
			12'b1101011011 		: log = 32'b00000000000000000011000010111101;
			12'b1101011100 		: log = 32'b00000000000000000011000011001010;
			12'b1101011101 		: log = 32'b00000000000000000011000011010111;
			12'b1101011110 		: log = 32'b00000000000000000011000011100100;
			12'b1101011111 		: log = 32'b00000000000000000011000011110010;
			12'b1101100000 		: log = 32'b00000000000000000011000011111111;
			12'b1101100001 		: log = 32'b00000000000000000011000100001100;
			12'b1101100010 		: log = 32'b00000000000000000011000100011001;
			12'b1101100011 		: log = 32'b00000000000000000011000100100110;
			12'b1101100100 		: log = 32'b00000000000000000011000100110100;
			12'b1101100101 		: log = 32'b00000000000000000011000101000001;
			12'b1101100110 		: log = 32'b00000000000000000011000101001110;
			12'b1101100111 		: log = 32'b00000000000000000011000101011011;
			12'b1101101000 		: log = 32'b00000000000000000011000101101000;
			12'b1101101001 		: log = 32'b00000000000000000011000101110110;
			12'b1101101010 		: log = 32'b00000000000000000011000110000011;
			12'b1101101011 		: log = 32'b00000000000000000011000110010000;
			12'b1101101100 		: log = 32'b00000000000000000011000110011101;
			12'b1101101101 		: log = 32'b00000000000000000011000110101010;
			12'b1101101110 		: log = 32'b00000000000000000011000110110111;
			12'b1101101111 		: log = 32'b00000000000000000011000111000101;
			12'b1101110000 		: log = 32'b00000000000000000011000111010010;
			12'b1101110001 		: log = 32'b00000000000000000011000111011111;
			12'b1101110010 		: log = 32'b00000000000000000011000111101100;
			12'b1101110011 		: log = 32'b00000000000000000011000111111001;
			12'b1101110100 		: log = 32'b00000000000000000011001000000110;
			12'b1101110101 		: log = 32'b00000000000000000011001000010100;
			12'b1101110110 		: log = 32'b00000000000000000011001000100001;
			12'b1101110111 		: log = 32'b00000000000000000011001000101110;
			12'b1101111000 		: log = 32'b00000000000000000011001000111011;
			12'b1101111001 		: log = 32'b00000000000000000011001001001000;
			12'b1101111010 		: log = 32'b00000000000000000011001001010101;
			12'b1101111011 		: log = 32'b00000000000000000011001001100011;
			12'b1101111100 		: log = 32'b00000000000000000011001001110000;
			12'b1101111101 		: log = 32'b00000000000000000011001001111101;
			12'b1101111110 		: log = 32'b00000000000000000011001010001010;
			12'b1101111111 		: log = 32'b00000000000000000011001010010111;
			12'b1110000000 		: log = 32'b00000000000000000011001010100100;
			12'b1110000001 		: log = 32'b00000000000000000011001010110001;
			12'b1110000010 		: log = 32'b00000000000000000011001010111110;
			12'b1110000011 		: log = 32'b00000000000000000011001011001100;
			12'b1110000100 		: log = 32'b00000000000000000011001011011001;
			12'b1110000101 		: log = 32'b00000000000000000011001011100110;
			12'b1110000110 		: log = 32'b00000000000000000011001011110011;
			12'b1110000111 		: log = 32'b00000000000000000011001100000000;
			12'b1110001000 		: log = 32'b00000000000000000011001100001101;
			12'b1110001001 		: log = 32'b00000000000000000011001100011010;
			12'b1110001010 		: log = 32'b00000000000000000011001100100111;
			12'b1110001011 		: log = 32'b00000000000000000011001100110100;
			12'b1110001100 		: log = 32'b00000000000000000011001101000010;
			12'b1110001101 		: log = 32'b00000000000000000011001101001111;
			12'b1110001110 		: log = 32'b00000000000000000011001101011100;
			12'b1110001111 		: log = 32'b00000000000000000011001101101001;
			12'b1110010000 		: log = 32'b00000000000000000011001101110110;
			12'b1110010001 		: log = 32'b00000000000000000011001110000011;
			12'b1110010010 		: log = 32'b00000000000000000011001110010000;
			12'b1110010011 		: log = 32'b00000000000000000011001110011101;
			12'b1110010100 		: log = 32'b00000000000000000011001110101010;
			12'b1110010101 		: log = 32'b00000000000000000011001110110111;
			12'b1110010110 		: log = 32'b00000000000000000011001111000100;
			12'b1110010111 		: log = 32'b00000000000000000011001111010001;
			12'b1110011000 		: log = 32'b00000000000000000011001111011111;
			12'b1110011001 		: log = 32'b00000000000000000011001111101100;
			12'b1110011010 		: log = 32'b00000000000000000011001111111001;
			12'b1110011011 		: log = 32'b00000000000000000011010000000110;
			12'b1110011100 		: log = 32'b00000000000000000011010000010011;
			12'b1110011101 		: log = 32'b00000000000000000011010000100000;
			12'b1110011110 		: log = 32'b00000000000000000011010000101101;
			12'b1110011111 		: log = 32'b00000000000000000011010000111010;
			12'b1110100000 		: log = 32'b00000000000000000011010001000111;
			12'b1110100001 		: log = 32'b00000000000000000011010001010100;
			12'b1110100010 		: log = 32'b00000000000000000011010001100001;
			12'b1110100011 		: log = 32'b00000000000000000011010001101110;
			12'b1110100100 		: log = 32'b00000000000000000011010001111011;
			12'b1110100101 		: log = 32'b00000000000000000011010010001000;
			12'b1110100110 		: log = 32'b00000000000000000011010010010101;
			12'b1110100111 		: log = 32'b00000000000000000011010010100010;
			12'b1110101000 		: log = 32'b00000000000000000011010010101111;
			12'b1110101001 		: log = 32'b00000000000000000011010010111100;
			12'b1110101010 		: log = 32'b00000000000000000011010011001001;
			12'b1110101011 		: log = 32'b00000000000000000011010011010110;
			12'b1110101100 		: log = 32'b00000000000000000011010011100011;
			12'b1110101101 		: log = 32'b00000000000000000011010011110000;
			12'b1110101110 		: log = 32'b00000000000000000011010011111101;
			12'b1110101111 		: log = 32'b00000000000000000011010100001010;
			12'b1110110000 		: log = 32'b00000000000000000011010100010111;
			12'b1110110001 		: log = 32'b00000000000000000011010100100100;
			12'b1110110010 		: log = 32'b00000000000000000011010100110001;
			12'b1110110011 		: log = 32'b00000000000000000011010100111110;
			12'b1110110100 		: log = 32'b00000000000000000011010101001011;
			12'b1110110101 		: log = 32'b00000000000000000011010101011000;
			12'b1110110110 		: log = 32'b00000000000000000011010101100101;
			12'b1110110111 		: log = 32'b00000000000000000011010101110010;
			12'b1110111000 		: log = 32'b00000000000000000011010101111111;
			12'b1110111001 		: log = 32'b00000000000000000011010110001100;
			12'b1110111010 		: log = 32'b00000000000000000011010110011001;
			12'b1110111011 		: log = 32'b00000000000000000011010110100110;
			12'b1110111100 		: log = 32'b00000000000000000011010110110011;
			12'b1110111101 		: log = 32'b00000000000000000011010111000000;
			12'b1110111110 		: log = 32'b00000000000000000011010111001101;
			12'b1110111111 		: log = 32'b00000000000000000011010111011010;
			12'b1111000000 		: log = 32'b00000000000000000011010111100111;
			12'b1111000001 		: log = 32'b00000000000000000011010111110100;
			12'b1111000010 		: log = 32'b00000000000000000011011000000001;
			12'b1111000011 		: log = 32'b00000000000000000011011000001110;
			12'b1111000100 		: log = 32'b00000000000000000011011000011011;
			12'b1111000101 		: log = 32'b00000000000000000011011000101000;
			12'b1111000110 		: log = 32'b00000000000000000011011000110101;
			12'b1111000111 		: log = 32'b00000000000000000011011001000010;
			12'b1111001000 		: log = 32'b00000000000000000011011001001111;
			12'b1111001001 		: log = 32'b00000000000000000011011001011100;
			12'b1111001010 		: log = 32'b00000000000000000011011001101001;
			12'b1111001011 		: log = 32'b00000000000000000011011001110110;
			12'b1111001100 		: log = 32'b00000000000000000011011010000010;
			12'b1111001101 		: log = 32'b00000000000000000011011010001111;
			12'b1111001110 		: log = 32'b00000000000000000011011010011100;
			12'b1111001111 		: log = 32'b00000000000000000011011010101001;
			12'b1111010000 		: log = 32'b00000000000000000011011010110110;
			12'b1111010001 		: log = 32'b00000000000000000011011011000011;
			12'b1111010010 		: log = 32'b00000000000000000011011011010000;
			12'b1111010011 		: log = 32'b00000000000000000011011011011101;
			12'b1111010100 		: log = 32'b00000000000000000011011011101010;
			12'b1111010101 		: log = 32'b00000000000000000011011011110111;
			12'b1111010110 		: log = 32'b00000000000000000011011100000100;
			12'b1111010111 		: log = 32'b00000000000000000011011100010001;
			12'b1111011000 		: log = 32'b00000000000000000011011100011101;
			12'b1111011001 		: log = 32'b00000000000000000011011100101010;
			12'b1111011010 		: log = 32'b00000000000000000011011100110111;
			12'b1111011011 		: log = 32'b00000000000000000011011101000100;
			12'b1111011100 		: log = 32'b00000000000000000011011101010001;
			12'b1111011101 		: log = 32'b00000000000000000011011101011110;
			12'b1111011110 		: log = 32'b00000000000000000011011101101011;
			12'b1111011111 		: log = 32'b00000000000000000011011101111000;
			12'b1111100000 		: log = 32'b00000000000000000011011110000101;
			12'b1111100001 		: log = 32'b00000000000000000011011110010001;
			12'b1111100010 		: log = 32'b00000000000000000011011110011110;
			12'b1111100011 		: log = 32'b00000000000000000011011110101011;
			12'b1111100100 		: log = 32'b00000000000000000011011110111000;
			12'b1111100101 		: log = 32'b00000000000000000011011111000101;
			12'b1111100110 		: log = 32'b00000000000000000011011111010010;
			12'b1111100111 		: log = 32'b00000000000000000011011111011111;
			12'b1111101000 		: log = 32'b00000000000000000011011111101100;
			12'b1111101001 		: log = 32'b00000000000000000011011111111000;
			12'b1111101010 		: log = 32'b00000000000000000011100000000101;
			12'b1111101011 		: log = 32'b00000000000000000011100000010010;
			12'b1111101100 		: log = 32'b00000000000000000011100000011111;
			12'b1111101101 		: log = 32'b00000000000000000011100000101100;
			12'b1111101110 		: log = 32'b00000000000000000011100000111001;
			12'b1111101111 		: log = 32'b00000000000000000011100001000101;
			12'b1111110000 		: log = 32'b00000000000000000011100001010010;
			12'b1111110001 		: log = 32'b00000000000000000011100001011111;
			12'b1111110010 		: log = 32'b00000000000000000011100001101100;
			12'b1111110011 		: log = 32'b00000000000000000011100001111001;
			12'b1111110100 		: log = 32'b00000000000000000011100010000110;
			12'b1111110101 		: log = 32'b00000000000000000011100010010010;
			12'b1111110110 		: log = 32'b00000000000000000011100010011111;
			12'b1111110111 		: log = 32'b00000000000000000011100010101100;
			12'b1111111000 		: log = 32'b00000000000000000011100010111001;
			12'b1111111001 		: log = 32'b00000000000000000011100011000110;
			12'b1111111010 		: log = 32'b00000000000000000011100011010011;
			12'b1111111011 		: log = 32'b00000000000000000011100011011111;
			12'b1111111100 		: log = 32'b00000000000000000011100011101100;
			12'b1111111101 		: log = 32'b00000000000000000011100011111001;
			12'b1111111110 		: log = 32'b00000000000000000011100100000110;
			12'b1111111111 		: log = 32'b00000000000000000011100100010011;
			12'b10000000000 		: log = 32'b00000000000000000011100100011111;
			12'b10000000001 		: log = 32'b00000000000000000011100100101100;
			12'b10000000010 		: log = 32'b00000000000000000011100100111001;
			12'b10000000011 		: log = 32'b00000000000000000011100101000110;
			12'b10000000100 		: log = 32'b00000000000000000011100101010011;
			12'b10000000101 		: log = 32'b00000000000000000011100101011111;
			12'b10000000110 		: log = 32'b00000000000000000011100101101100;
			12'b10000000111 		: log = 32'b00000000000000000011100101111001;
			12'b10000001000 		: log = 32'b00000000000000000011100110000110;
			12'b10000001001 		: log = 32'b00000000000000000011100110010011;
			12'b10000001010 		: log = 32'b00000000000000000011100110011111;
			12'b10000001011 		: log = 32'b00000000000000000011100110101100;
			12'b10000001100 		: log = 32'b00000000000000000011100110111001;
			12'b10000001101 		: log = 32'b00000000000000000011100111000110;
			12'b10000001110 		: log = 32'b00000000000000000011100111010010;
			12'b10000001111 		: log = 32'b00000000000000000011100111011111;
			12'b10000010000 		: log = 32'b00000000000000000011100111101100;
			12'b10000010001 		: log = 32'b00000000000000000011100111111001;
			12'b10000010010 		: log = 32'b00000000000000000011101000000101;
			12'b10000010011 		: log = 32'b00000000000000000011101000010010;
			12'b10000010100 		: log = 32'b00000000000000000011101000011111;
			12'b10000010101 		: log = 32'b00000000000000000011101000101100;
			12'b10000010110 		: log = 32'b00000000000000000011101000111000;
			12'b10000010111 		: log = 32'b00000000000000000011101001000101;
			12'b10000011000 		: log = 32'b00000000000000000011101001010010;
			12'b10000011001 		: log = 32'b00000000000000000011101001011111;
			12'b10000011010 		: log = 32'b00000000000000000011101001101011;
			12'b10000011011 		: log = 32'b00000000000000000011101001111000;
			12'b10000011100 		: log = 32'b00000000000000000011101010000101;
			12'b10000011101 		: log = 32'b00000000000000000011101010010010;
			12'b10000011110 		: log = 32'b00000000000000000011101010011110;
			12'b10000011111 		: log = 32'b00000000000000000011101010101011;
			12'b10000100000 		: log = 32'b00000000000000000011101010111000;
			12'b10000100001 		: log = 32'b00000000000000000011101011000100;
			12'b10000100010 		: log = 32'b00000000000000000011101011010001;
			12'b10000100011 		: log = 32'b00000000000000000011101011011110;
			12'b10000100100 		: log = 32'b00000000000000000011101011101011;
			12'b10000100101 		: log = 32'b00000000000000000011101011110111;
			12'b10000100110 		: log = 32'b00000000000000000011101100000100;
			12'b10000100111 		: log = 32'b00000000000000000011101100010001;
			12'b10000101000 		: log = 32'b00000000000000000011101100011101;
			12'b10000101001 		: log = 32'b00000000000000000011101100101010;
			12'b10000101010 		: log = 32'b00000000000000000011101100110111;
			12'b10000101011 		: log = 32'b00000000000000000011101101000100;
			12'b10000101100 		: log = 32'b00000000000000000011101101010000;
			12'b10000101101 		: log = 32'b00000000000000000011101101011101;
			12'b10000101110 		: log = 32'b00000000000000000011101101101010;
			12'b10000101111 		: log = 32'b00000000000000000011101101110110;
			12'b10000110000 		: log = 32'b00000000000000000011101110000011;
			12'b10000110001 		: log = 32'b00000000000000000011101110010000;
			12'b10000110010 		: log = 32'b00000000000000000011101110011100;
			12'b10000110011 		: log = 32'b00000000000000000011101110101001;
			12'b10000110100 		: log = 32'b00000000000000000011101110110110;
			12'b10000110101 		: log = 32'b00000000000000000011101111000010;
			12'b10000110110 		: log = 32'b00000000000000000011101111001111;
			12'b10000110111 		: log = 32'b00000000000000000011101111011100;
			12'b10000111000 		: log = 32'b00000000000000000011101111101000;
			12'b10000111001 		: log = 32'b00000000000000000011101111110101;
			12'b10000111010 		: log = 32'b00000000000000000011110000000010;
			12'b10000111011 		: log = 32'b00000000000000000011110000001110;
			12'b10000111100 		: log = 32'b00000000000000000011110000011011;
			12'b10000111101 		: log = 32'b00000000000000000011110000101000;
			12'b10000111110 		: log = 32'b00000000000000000011110000110100;
			12'b10000111111 		: log = 32'b00000000000000000011110001000001;
			12'b10001000000 		: log = 32'b00000000000000000011110001001110;
			12'b10001000001 		: log = 32'b00000000000000000011110001011010;
			12'b10001000010 		: log = 32'b00000000000000000011110001100111;
			12'b10001000011 		: log = 32'b00000000000000000011110001110011;
			12'b10001000100 		: log = 32'b00000000000000000011110010000000;
			12'b10001000101 		: log = 32'b00000000000000000011110010001101;
			12'b10001000110 		: log = 32'b00000000000000000011110010011001;
			12'b10001000111 		: log = 32'b00000000000000000011110010100110;
			12'b10001001000 		: log = 32'b00000000000000000011110010110011;
			12'b10001001001 		: log = 32'b00000000000000000011110010111111;
			12'b10001001010 		: log = 32'b00000000000000000011110011001100;
			12'b10001001011 		: log = 32'b00000000000000000011110011011000;
			12'b10001001100 		: log = 32'b00000000000000000011110011100101;
			12'b10001001101 		: log = 32'b00000000000000000011110011110010;
			12'b10001001110 		: log = 32'b00000000000000000011110011111110;
			12'b10001001111 		: log = 32'b00000000000000000011110100001011;
			12'b10001010000 		: log = 32'b00000000000000000011110100011000;
			12'b10001010001 		: log = 32'b00000000000000000011110100100100;
			12'b10001010010 		: log = 32'b00000000000000000011110100110001;
			12'b10001010011 		: log = 32'b00000000000000000011110100111101;
			12'b10001010100 		: log = 32'b00000000000000000011110101001010;
			12'b10001010101 		: log = 32'b00000000000000000011110101010111;
			12'b10001010110 		: log = 32'b00000000000000000011110101100011;
			12'b10001010111 		: log = 32'b00000000000000000011110101110000;
			12'b10001011000 		: log = 32'b00000000000000000011110101111100;
			12'b10001011001 		: log = 32'b00000000000000000011110110001001;
			12'b10001011010 		: log = 32'b00000000000000000011110110010101;
			12'b10001011011 		: log = 32'b00000000000000000011110110100010;
			12'b10001011100 		: log = 32'b00000000000000000011110110101111;
			12'b10001011101 		: log = 32'b00000000000000000011110110111011;
			12'b10001011110 		: log = 32'b00000000000000000011110111001000;
			12'b10001011111 		: log = 32'b00000000000000000011110111010100;
			12'b10001100000 		: log = 32'b00000000000000000011110111100001;
			12'b10001100001 		: log = 32'b00000000000000000011110111101101;
			12'b10001100010 		: log = 32'b00000000000000000011110111111010;
			12'b10001100011 		: log = 32'b00000000000000000011111000000111;
			12'b10001100100 		: log = 32'b00000000000000000011111000010011;
			12'b10001100101 		: log = 32'b00000000000000000011111000100000;
			12'b10001100110 		: log = 32'b00000000000000000011111000101100;
			12'b10001100111 		: log = 32'b00000000000000000011111000111001;
			12'b10001101000 		: log = 32'b00000000000000000011111001000101;
			12'b10001101001 		: log = 32'b00000000000000000011111001010010;
			12'b10001101010 		: log = 32'b00000000000000000011111001011110;
			12'b10001101011 		: log = 32'b00000000000000000011111001101011;
			12'b10001101100 		: log = 32'b00000000000000000011111001110111;
			12'b10001101101 		: log = 32'b00000000000000000011111010000100;
			12'b10001101110 		: log = 32'b00000000000000000011111010010001;
			12'b10001101111 		: log = 32'b00000000000000000011111010011101;
			12'b10001110000 		: log = 32'b00000000000000000011111010101010;
			12'b10001110001 		: log = 32'b00000000000000000011111010110110;
			12'b10001110010 		: log = 32'b00000000000000000011111011000011;
			12'b10001110011 		: log = 32'b00000000000000000011111011001111;
			12'b10001110100 		: log = 32'b00000000000000000011111011011100;
			12'b10001110101 		: log = 32'b00000000000000000011111011101000;
			12'b10001110110 		: log = 32'b00000000000000000011111011110101;
			12'b10001110111 		: log = 32'b00000000000000000011111100000001;
			12'b10001111000 		: log = 32'b00000000000000000011111100001110;
			12'b10001111001 		: log = 32'b00000000000000000011111100011010;
			12'b10001111010 		: log = 32'b00000000000000000011111100100111;
			12'b10001111011 		: log = 32'b00000000000000000011111100110011;
			12'b10001111100 		: log = 32'b00000000000000000011111101000000;
			12'b10001111101 		: log = 32'b00000000000000000011111101001100;
			12'b10001111110 		: log = 32'b00000000000000000011111101011001;
			12'b10001111111 		: log = 32'b00000000000000000011111101100101;
			12'b10010000000 		: log = 32'b00000000000000000011111101110010;
			12'b10010000001 		: log = 32'b00000000000000000011111101111110;
			12'b10010000010 		: log = 32'b00000000000000000011111110001011;
			12'b10010000011 		: log = 32'b00000000000000000011111110010111;
			12'b10010000100 		: log = 32'b00000000000000000011111110100100;
			12'b10010000101 		: log = 32'b00000000000000000011111110110000;
			12'b10010000110 		: log = 32'b00000000000000000011111110111101;
			12'b10010000111 		: log = 32'b00000000000000000011111111001001;
			12'b10010001000 		: log = 32'b00000000000000000011111111010110;
			12'b10010001001 		: log = 32'b00000000000000000011111111100010;
			12'b10010001010 		: log = 32'b00000000000000000011111111101110;
			12'b10010001011 		: log = 32'b00000000000000000011111111111011;
			12'b10010001100 		: log = 32'b00000000000000000100000000000111;
			12'b10010001101 		: log = 32'b00000000000000000100000000010100;
			12'b10010001110 		: log = 32'b00000000000000000100000000100000;
			12'b10010001111 		: log = 32'b00000000000000000100000000101101;
			12'b10010010000 		: log = 32'b00000000000000000100000000111001;
			12'b10010010001 		: log = 32'b00000000000000000100000001000110;
			12'b10010010010 		: log = 32'b00000000000000000100000001010010;
			12'b10010010011 		: log = 32'b00000000000000000100000001011111;
			12'b10010010100 		: log = 32'b00000000000000000100000001101011;
			12'b10010010101 		: log = 32'b00000000000000000100000001110111;
			12'b10010010110 		: log = 32'b00000000000000000100000010000100;
			12'b10010010111 		: log = 32'b00000000000000000100000010010000;
			12'b10010011000 		: log = 32'b00000000000000000100000010011101;
			12'b10010011001 		: log = 32'b00000000000000000100000010101001;
			12'b10010011010 		: log = 32'b00000000000000000100000010110110;
			12'b10010011011 		: log = 32'b00000000000000000100000011000010;
			12'b10010011100 		: log = 32'b00000000000000000100000011001110;
			12'b10010011101 		: log = 32'b00000000000000000100000011011011;
			12'b10010011110 		: log = 32'b00000000000000000100000011100111;
			12'b10010011111 		: log = 32'b00000000000000000100000011110100;
			12'b10010100000 		: log = 32'b00000000000000000100000100000000;
			12'b10010100001 		: log = 32'b00000000000000000100000100001100;
			12'b10010100010 		: log = 32'b00000000000000000100000100011001;
			12'b10010100011 		: log = 32'b00000000000000000100000100100101;
			12'b10010100100 		: log = 32'b00000000000000000100000100110010;
			12'b10010100101 		: log = 32'b00000000000000000100000100111110;
			12'b10010100110 		: log = 32'b00000000000000000100000101001011;
			12'b10010100111 		: log = 32'b00000000000000000100000101010111;
			12'b10010101000 		: log = 32'b00000000000000000100000101100011;
			12'b10010101001 		: log = 32'b00000000000000000100000101110000;
			12'b10010101010 		: log = 32'b00000000000000000100000101111100;
			12'b10010101011 		: log = 32'b00000000000000000100000110001000;
			12'b10010101100 		: log = 32'b00000000000000000100000110010101;
			12'b10010101101 		: log = 32'b00000000000000000100000110100001;
			12'b10010101110 		: log = 32'b00000000000000000100000110101110;
			12'b10010101111 		: log = 32'b00000000000000000100000110111010;
			12'b10010110000 		: log = 32'b00000000000000000100000111000110;
			12'b10010110001 		: log = 32'b00000000000000000100000111010011;
			12'b10010110010 		: log = 32'b00000000000000000100000111011111;
			12'b10010110011 		: log = 32'b00000000000000000100000111101011;
			12'b10010110100 		: log = 32'b00000000000000000100000111111000;
			12'b10010110101 		: log = 32'b00000000000000000100001000000100;
			12'b10010110110 		: log = 32'b00000000000000000100001000010001;
			12'b10010110111 		: log = 32'b00000000000000000100001000011101;
			12'b10010111000 		: log = 32'b00000000000000000100001000101001;
			12'b10010111001 		: log = 32'b00000000000000000100001000110110;
			12'b10010111010 		: log = 32'b00000000000000000100001001000010;
			12'b10010111011 		: log = 32'b00000000000000000100001001001110;
			12'b10010111100 		: log = 32'b00000000000000000100001001011011;
			12'b10010111101 		: log = 32'b00000000000000000100001001100111;
			12'b10010111110 		: log = 32'b00000000000000000100001001110011;
			12'b10010111111 		: log = 32'b00000000000000000100001010000000;
			12'b10011000000 		: log = 32'b00000000000000000100001010001100;
			12'b10011000001 		: log = 32'b00000000000000000100001010011000;
			12'b10011000010 		: log = 32'b00000000000000000100001010100101;
			12'b10011000011 		: log = 32'b00000000000000000100001010110001;
			12'b10011000100 		: log = 32'b00000000000000000100001010111101;
			12'b10011000101 		: log = 32'b00000000000000000100001011001010;
			12'b10011000110 		: log = 32'b00000000000000000100001011010110;
			12'b10011000111 		: log = 32'b00000000000000000100001011100010;
			12'b10011001000 		: log = 32'b00000000000000000100001011101111;
			12'b10011001001 		: log = 32'b00000000000000000100001011111011;
			12'b10011001010 		: log = 32'b00000000000000000100001100000111;
			12'b10011001011 		: log = 32'b00000000000000000100001100010100;
			12'b10011001100 		: log = 32'b00000000000000000100001100100000;
			12'b10011001101 		: log = 32'b00000000000000000100001100101100;
			12'b10011001110 		: log = 32'b00000000000000000100001100111001;
			12'b10011001111 		: log = 32'b00000000000000000100001101000101;
			12'b10011010000 		: log = 32'b00000000000000000100001101010001;
			12'b10011010001 		: log = 32'b00000000000000000100001101011101;
			12'b10011010010 		: log = 32'b00000000000000000100001101101010;
			12'b10011010011 		: log = 32'b00000000000000000100001101110110;
			12'b10011010100 		: log = 32'b00000000000000000100001110000010;
			12'b10011010101 		: log = 32'b00000000000000000100001110001111;
			12'b10011010110 		: log = 32'b00000000000000000100001110011011;
			12'b10011010111 		: log = 32'b00000000000000000100001110100111;
			12'b10011011000 		: log = 32'b00000000000000000100001110110100;
			12'b10011011001 		: log = 32'b00000000000000000100001111000000;
			12'b10011011010 		: log = 32'b00000000000000000100001111001100;
			12'b10011011011 		: log = 32'b00000000000000000100001111011000;
			12'b10011011100 		: log = 32'b00000000000000000100001111100101;
			12'b10011011101 		: log = 32'b00000000000000000100001111110001;
			12'b10011011110 		: log = 32'b00000000000000000100001111111101;
			12'b10011011111 		: log = 32'b00000000000000000100010000001001;
			12'b10011100000 		: log = 32'b00000000000000000100010000010110;
			12'b10011100001 		: log = 32'b00000000000000000100010000100010;
			12'b10011100010 		: log = 32'b00000000000000000100010000101110;
			12'b10011100011 		: log = 32'b00000000000000000100010000111010;
			12'b10011100100 		: log = 32'b00000000000000000100010001000111;
			12'b10011100101 		: log = 32'b00000000000000000100010001010011;
			12'b10011100110 		: log = 32'b00000000000000000100010001011111;
			12'b10011100111 		: log = 32'b00000000000000000100010001101011;
			12'b10011101000 		: log = 32'b00000000000000000100010001111000;
			12'b10011101001 		: log = 32'b00000000000000000100010010000100;
			12'b10011101010 		: log = 32'b00000000000000000100010010010000;
			12'b10011101011 		: log = 32'b00000000000000000100010010011100;
			12'b10011101100 		: log = 32'b00000000000000000100010010101001;
			12'b10011101101 		: log = 32'b00000000000000000100010010110101;
			12'b10011101110 		: log = 32'b00000000000000000100010011000001;
			12'b10011101111 		: log = 32'b00000000000000000100010011001101;
			12'b10011110000 		: log = 32'b00000000000000000100010011011010;
			12'b10011110001 		: log = 32'b00000000000000000100010011100110;
			12'b10011110010 		: log = 32'b00000000000000000100010011110010;
			12'b10011110011 		: log = 32'b00000000000000000100010011111110;
			12'b10011110100 		: log = 32'b00000000000000000100010100001010;
			12'b10011110101 		: log = 32'b00000000000000000100010100010111;
			12'b10011110110 		: log = 32'b00000000000000000100010100100011;
			12'b10011110111 		: log = 32'b00000000000000000100010100101111;
			12'b10011111000 		: log = 32'b00000000000000000100010100111011;
			12'b10011111001 		: log = 32'b00000000000000000100010101001000;
			12'b10011111010 		: log = 32'b00000000000000000100010101010100;
			12'b10011111011 		: log = 32'b00000000000000000100010101100000;
			12'b10011111100 		: log = 32'b00000000000000000100010101101100;
			12'b10011111101 		: log = 32'b00000000000000000100010101111000;
			12'b10011111110 		: log = 32'b00000000000000000100010110000101;
			12'b10011111111 		: log = 32'b00000000000000000100010110010001;
			12'b10100000000 		: log = 32'b00000000000000000100010110011101;
			12'b10100000001 		: log = 32'b00000000000000000100010110101001;
			12'b10100000010 		: log = 32'b00000000000000000100010110110101;
			12'b10100000011 		: log = 32'b00000000000000000100010111000010;
			12'b10100000100 		: log = 32'b00000000000000000100010111001110;
			12'b10100000101 		: log = 32'b00000000000000000100010111011010;
			12'b10100000110 		: log = 32'b00000000000000000100010111100110;
			12'b10100000111 		: log = 32'b00000000000000000100010111110010;
			12'b10100001000 		: log = 32'b00000000000000000100010111111110;
			12'b10100001001 		: log = 32'b00000000000000000100011000001011;
			12'b10100001010 		: log = 32'b00000000000000000100011000010111;
			12'b10100001011 		: log = 32'b00000000000000000100011000100011;
			12'b10100001100 		: log = 32'b00000000000000000100011000101111;
			12'b10100001101 		: log = 32'b00000000000000000100011000111011;
			12'b10100001110 		: log = 32'b00000000000000000100011001000111;
			12'b10100001111 		: log = 32'b00000000000000000100011001010100;
			12'b10100010000 		: log = 32'b00000000000000000100011001100000;
			12'b10100010001 		: log = 32'b00000000000000000100011001101100;
			12'b10100010010 		: log = 32'b00000000000000000100011001111000;
			12'b10100010011 		: log = 32'b00000000000000000100011010000100;
			12'b10100010100 		: log = 32'b00000000000000000100011010010000;
			12'b10100010101 		: log = 32'b00000000000000000100011010011100;
			12'b10100010110 		: log = 32'b00000000000000000100011010101001;
			12'b10100010111 		: log = 32'b00000000000000000100011010110101;
			12'b10100011000 		: log = 32'b00000000000000000100011011000001;
			12'b10100011001 		: log = 32'b00000000000000000100011011001101;
			12'b10100011010 		: log = 32'b00000000000000000100011011011001;
			12'b10100011011 		: log = 32'b00000000000000000100011011100101;
			12'b10100011100 		: log = 32'b00000000000000000100011011110001;
			12'b10100011101 		: log = 32'b00000000000000000100011011111110;
			12'b10100011110 		: log = 32'b00000000000000000100011100001010;
			12'b10100011111 		: log = 32'b00000000000000000100011100010110;
			12'b10100100000 		: log = 32'b00000000000000000100011100100010;
			12'b10100100001 		: log = 32'b00000000000000000100011100101110;
			12'b10100100010 		: log = 32'b00000000000000000100011100111010;
			12'b10100100011 		: log = 32'b00000000000000000100011101000110;
			12'b10100100100 		: log = 32'b00000000000000000100011101010010;
			12'b10100100101 		: log = 32'b00000000000000000100011101011110;
			12'b10100100110 		: log = 32'b00000000000000000100011101101011;
			12'b10100100111 		: log = 32'b00000000000000000100011101110111;
			12'b10100101000 		: log = 32'b00000000000000000100011110000011;
			12'b10100101001 		: log = 32'b00000000000000000100011110001111;
			12'b10100101010 		: log = 32'b00000000000000000100011110011011;
			12'b10100101011 		: log = 32'b00000000000000000100011110100111;
			12'b10100101100 		: log = 32'b00000000000000000100011110110011;
			12'b10100101101 		: log = 32'b00000000000000000100011110111111;
			12'b10100101110 		: log = 32'b00000000000000000100011111001011;
			12'b10100101111 		: log = 32'b00000000000000000100011111010111;
			12'b10100110000 		: log = 32'b00000000000000000100011111100011;
			12'b10100110001 		: log = 32'b00000000000000000100011111110000;
			12'b10100110010 		: log = 32'b00000000000000000100011111111100;
			12'b10100110011 		: log = 32'b00000000000000000100100000001000;
			12'b10100110100 		: log = 32'b00000000000000000100100000010100;
			12'b10100110101 		: log = 32'b00000000000000000100100000100000;
			12'b10100110110 		: log = 32'b00000000000000000100100000101100;
			12'b10100110111 		: log = 32'b00000000000000000100100000111000;
			12'b10100111000 		: log = 32'b00000000000000000100100001000100;
			12'b10100111001 		: log = 32'b00000000000000000100100001010000;
			12'b10100111010 		: log = 32'b00000000000000000100100001011100;
			12'b10100111011 		: log = 32'b00000000000000000100100001101000;
			12'b10100111100 		: log = 32'b00000000000000000100100001110100;
			12'b10100111101 		: log = 32'b00000000000000000100100010000000;
			12'b10100111110 		: log = 32'b00000000000000000100100010001100;
			12'b10100111111 		: log = 32'b00000000000000000100100010011000;
			12'b10101000000 		: log = 32'b00000000000000000100100010100101;
			12'b10101000001 		: log = 32'b00000000000000000100100010110001;
			12'b10101000010 		: log = 32'b00000000000000000100100010111101;
			12'b10101000011 		: log = 32'b00000000000000000100100011001001;
			12'b10101000100 		: log = 32'b00000000000000000100100011010101;
			12'b10101000101 		: log = 32'b00000000000000000100100011100001;
			12'b10101000110 		: log = 32'b00000000000000000100100011101101;
			12'b10101000111 		: log = 32'b00000000000000000100100011111001;
			12'b10101001000 		: log = 32'b00000000000000000100100100000101;
			12'b10101001001 		: log = 32'b00000000000000000100100100010001;
			12'b10101001010 		: log = 32'b00000000000000000100100100011101;
			12'b10101001011 		: log = 32'b00000000000000000100100100101001;
			12'b10101001100 		: log = 32'b00000000000000000100100100110101;
			12'b10101001101 		: log = 32'b00000000000000000100100101000001;
			12'b10101001110 		: log = 32'b00000000000000000100100101001101;
			12'b10101001111 		: log = 32'b00000000000000000100100101011001;
			12'b10101010000 		: log = 32'b00000000000000000100100101100101;
			12'b10101010001 		: log = 32'b00000000000000000100100101110001;
			12'b10101010010 		: log = 32'b00000000000000000100100101111101;
			12'b10101010011 		: log = 32'b00000000000000000100100110001001;
			12'b10101010100 		: log = 32'b00000000000000000100100110010101;
			12'b10101010101 		: log = 32'b00000000000000000100100110100001;
			12'b10101010110 		: log = 32'b00000000000000000100100110101101;
			12'b10101010111 		: log = 32'b00000000000000000100100110111001;
			12'b10101011000 		: log = 32'b00000000000000000100100111000101;
			12'b10101011001 		: log = 32'b00000000000000000100100111010001;
			12'b10101011010 		: log = 32'b00000000000000000100100111011101;
			12'b10101011011 		: log = 32'b00000000000000000100100111101001;
			12'b10101011100 		: log = 32'b00000000000000000100100111110101;
			12'b10101011101 		: log = 32'b00000000000000000100101000000001;
			12'b10101011110 		: log = 32'b00000000000000000100101000001101;
			12'b10101011111 		: log = 32'b00000000000000000100101000011001;
			12'b10101100000 		: log = 32'b00000000000000000100101000100101;
			12'b10101100001 		: log = 32'b00000000000000000100101000110001;
			12'b10101100010 		: log = 32'b00000000000000000100101000111101;
			12'b10101100011 		: log = 32'b00000000000000000100101001001001;
			12'b10101100100 		: log = 32'b00000000000000000100101001010101;
			12'b10101100101 		: log = 32'b00000000000000000100101001100001;
			12'b10101100110 		: log = 32'b00000000000000000100101001101101;
			12'b10101100111 		: log = 32'b00000000000000000100101001111001;
			12'b10101101000 		: log = 32'b00000000000000000100101010000101;
			12'b10101101001 		: log = 32'b00000000000000000100101010010001;
			12'b10101101010 		: log = 32'b00000000000000000100101010011101;
			12'b10101101011 		: log = 32'b00000000000000000100101010101001;
			12'b10101101100 		: log = 32'b00000000000000000100101010110100;
			12'b10101101101 		: log = 32'b00000000000000000100101011000000;
			12'b10101101110 		: log = 32'b00000000000000000100101011001100;
			12'b10101101111 		: log = 32'b00000000000000000100101011011000;
			12'b10101110000 		: log = 32'b00000000000000000100101011100100;
			12'b10101110001 		: log = 32'b00000000000000000100101011110000;
			12'b10101110010 		: log = 32'b00000000000000000100101011111100;
			12'b10101110011 		: log = 32'b00000000000000000100101100001000;
			12'b10101110100 		: log = 32'b00000000000000000100101100010100;
			12'b10101110101 		: log = 32'b00000000000000000100101100100000;
			12'b10101110110 		: log = 32'b00000000000000000100101100101100;
			12'b10101110111 		: log = 32'b00000000000000000100101100111000;
			12'b10101111000 		: log = 32'b00000000000000000100101101000100;
			12'b10101111001 		: log = 32'b00000000000000000100101101010000;
			12'b10101111010 		: log = 32'b00000000000000000100101101011100;
			12'b10101111011 		: log = 32'b00000000000000000100101101100111;
			12'b10101111100 		: log = 32'b00000000000000000100101101110011;
			12'b10101111101 		: log = 32'b00000000000000000100101101111111;
			12'b10101111110 		: log = 32'b00000000000000000100101110001011;
			12'b10101111111 		: log = 32'b00000000000000000100101110010111;
			12'b10110000000 		: log = 32'b00000000000000000100101110100011;
			12'b10110000001 		: log = 32'b00000000000000000100101110101111;
			12'b10110000010 		: log = 32'b00000000000000000100101110111011;
			12'b10110000011 		: log = 32'b00000000000000000100101111000111;
			12'b10110000100 		: log = 32'b00000000000000000100101111010011;
			12'b10110000101 		: log = 32'b00000000000000000100101111011111;
			12'b10110000110 		: log = 32'b00000000000000000100101111101010;
			12'b10110000111 		: log = 32'b00000000000000000100101111110110;
			12'b10110001000 		: log = 32'b00000000000000000100110000000010;
			12'b10110001001 		: log = 32'b00000000000000000100110000001110;
			12'b10110001010 		: log = 32'b00000000000000000100110000011010;
			12'b10110001011 		: log = 32'b00000000000000000100110000100110;
			12'b10110001100 		: log = 32'b00000000000000000100110000110010;
			12'b10110001101 		: log = 32'b00000000000000000100110000111110;
			12'b10110001110 		: log = 32'b00000000000000000100110001001010;
			12'b10110001111 		: log = 32'b00000000000000000100110001010101;
			12'b10110010000 		: log = 32'b00000000000000000100110001100001;
			12'b10110010001 		: log = 32'b00000000000000000100110001101101;
			12'b10110010010 		: log = 32'b00000000000000000100110001111001;
			12'b10110010011 		: log = 32'b00000000000000000100110010000101;
			12'b10110010100 		: log = 32'b00000000000000000100110010010001;
			12'b10110010101 		: log = 32'b00000000000000000100110010011101;
			12'b10110010110 		: log = 32'b00000000000000000100110010101000;
			12'b10110010111 		: log = 32'b00000000000000000100110010110100;
			12'b10110011000 		: log = 32'b00000000000000000100110011000000;
			12'b10110011001 		: log = 32'b00000000000000000100110011001100;
			12'b10110011010 		: log = 32'b00000000000000000100110011011000;
			12'b10110011011 		: log = 32'b00000000000000000100110011100100;
			12'b10110011100 		: log = 32'b00000000000000000100110011110000;
			12'b10110011101 		: log = 32'b00000000000000000100110011111011;
			12'b10110011110 		: log = 32'b00000000000000000100110100000111;
			12'b10110011111 		: log = 32'b00000000000000000100110100010011;
			12'b10110100000 		: log = 32'b00000000000000000100110100011111;
			12'b10110100001 		: log = 32'b00000000000000000100110100101011;
			12'b10110100010 		: log = 32'b00000000000000000100110100110111;
			12'b10110100011 		: log = 32'b00000000000000000100110101000010;
			12'b10110100100 		: log = 32'b00000000000000000100110101001110;
			12'b10110100101 		: log = 32'b00000000000000000100110101011010;
			12'b10110100110 		: log = 32'b00000000000000000100110101100110;
			12'b10110100111 		: log = 32'b00000000000000000100110101110010;
			12'b10110101000 		: log = 32'b00000000000000000100110101111110;
			12'b10110101001 		: log = 32'b00000000000000000100110110001001;
			12'b10110101010 		: log = 32'b00000000000000000100110110010101;
			12'b10110101011 		: log = 32'b00000000000000000100110110100001;
			12'b10110101100 		: log = 32'b00000000000000000100110110101101;
			12'b10110101101 		: log = 32'b00000000000000000100110110111001;
			12'b10110101110 		: log = 32'b00000000000000000100110111000100;
			12'b10110101111 		: log = 32'b00000000000000000100110111010000;
			12'b10110110000 		: log = 32'b00000000000000000100110111011100;
			12'b10110110001 		: log = 32'b00000000000000000100110111101000;
			12'b10110110010 		: log = 32'b00000000000000000100110111110100;
			12'b10110110011 		: log = 32'b00000000000000000100111000000000;
			12'b10110110100 		: log = 32'b00000000000000000100111000001011;
			12'b10110110101 		: log = 32'b00000000000000000100111000010111;
			12'b10110110110 		: log = 32'b00000000000000000100111000100011;
			12'b10110110111 		: log = 32'b00000000000000000100111000101111;
			12'b10110111000 		: log = 32'b00000000000000000100111000111010;
			12'b10110111001 		: log = 32'b00000000000000000100111001000110;
			12'b10110111010 		: log = 32'b00000000000000000100111001010010;
			12'b10110111011 		: log = 32'b00000000000000000100111001011110;
			12'b10110111100 		: log = 32'b00000000000000000100111001101010;
			12'b10110111101 		: log = 32'b00000000000000000100111001110101;
			12'b10110111110 		: log = 32'b00000000000000000100111010000001;
			12'b10110111111 		: log = 32'b00000000000000000100111010001101;
			12'b10111000000 		: log = 32'b00000000000000000100111010011001;
			12'b10111000001 		: log = 32'b00000000000000000100111010100100;
			12'b10111000010 		: log = 32'b00000000000000000100111010110000;
			12'b10111000011 		: log = 32'b00000000000000000100111010111100;
			12'b10111000100 		: log = 32'b00000000000000000100111011001000;
			12'b10111000101 		: log = 32'b00000000000000000100111011010100;
			12'b10111000110 		: log = 32'b00000000000000000100111011011111;
			12'b10111000111 		: log = 32'b00000000000000000100111011101011;
			12'b10111001000 		: log = 32'b00000000000000000100111011110111;
			12'b10111001001 		: log = 32'b00000000000000000100111100000011;
			12'b10111001010 		: log = 32'b00000000000000000100111100001110;
			12'b10111001011 		: log = 32'b00000000000000000100111100011010;
			12'b10111001100 		: log = 32'b00000000000000000100111100100110;
			12'b10111001101 		: log = 32'b00000000000000000100111100110010;
			12'b10111001110 		: log = 32'b00000000000000000100111100111101;
			12'b10111001111 		: log = 32'b00000000000000000100111101001001;
			12'b10111010000 		: log = 32'b00000000000000000100111101010101;
			12'b10111010001 		: log = 32'b00000000000000000100111101100000;
			12'b10111010010 		: log = 32'b00000000000000000100111101101100;
			12'b10111010011 		: log = 32'b00000000000000000100111101111000;
			12'b10111010100 		: log = 32'b00000000000000000100111110000100;
			12'b10111010101 		: log = 32'b00000000000000000100111110001111;
			12'b10111010110 		: log = 32'b00000000000000000100111110011011;
			12'b10111010111 		: log = 32'b00000000000000000100111110100111;
			12'b10111011000 		: log = 32'b00000000000000000100111110110011;
			12'b10111011001 		: log = 32'b00000000000000000100111110111110;
			12'b10111011010 		: log = 32'b00000000000000000100111111001010;
			12'b10111011011 		: log = 32'b00000000000000000100111111010110;
			12'b10111011100 		: log = 32'b00000000000000000100111111100001;
			12'b10111011101 		: log = 32'b00000000000000000100111111101101;
			12'b10111011110 		: log = 32'b00000000000000000100111111111001;
			12'b10111011111 		: log = 32'b00000000000000000101000000000101;
			12'b10111100000 		: log = 32'b00000000000000000101000000010000;
			12'b10111100001 		: log = 32'b00000000000000000101000000011100;
			12'b10111100010 		: log = 32'b00000000000000000101000000101000;
			12'b10111100011 		: log = 32'b00000000000000000101000000110011;
			12'b10111100100 		: log = 32'b00000000000000000101000000111111;
			12'b10111100101 		: log = 32'b00000000000000000101000001001011;
			12'b10111100110 		: log = 32'b00000000000000000101000001010110;
			12'b10111100111 		: log = 32'b00000000000000000101000001100010;
			12'b10111101000 		: log = 32'b00000000000000000101000001101110;
			12'b10111101001 		: log = 32'b00000000000000000101000001111001;
			12'b10111101010 		: log = 32'b00000000000000000101000010000101;
			12'b10111101011 		: log = 32'b00000000000000000101000010010001;
			12'b10111101100 		: log = 32'b00000000000000000101000010011101;
			12'b10111101101 		: log = 32'b00000000000000000101000010101000;
			12'b10111101110 		: log = 32'b00000000000000000101000010110100;
			12'b10111101111 		: log = 32'b00000000000000000101000011000000;
			12'b10111110000 		: log = 32'b00000000000000000101000011001011;
			12'b10111110001 		: log = 32'b00000000000000000101000011010111;
			12'b10111110010 		: log = 32'b00000000000000000101000011100011;
			12'b10111110011 		: log = 32'b00000000000000000101000011101110;
			12'b10111110100 		: log = 32'b00000000000000000101000011111010;
			12'b10111110101 		: log = 32'b00000000000000000101000100000110;
			12'b10111110110 		: log = 32'b00000000000000000101000100010001;
			12'b10111110111 		: log = 32'b00000000000000000101000100011101;
			12'b10111111000 		: log = 32'b00000000000000000101000100101001;
			12'b10111111001 		: log = 32'b00000000000000000101000100110100;
			12'b10111111010 		: log = 32'b00000000000000000101000101000000;
			12'b10111111011 		: log = 32'b00000000000000000101000101001011;
			12'b10111111100 		: log = 32'b00000000000000000101000101010111;
			12'b10111111101 		: log = 32'b00000000000000000101000101100011;
			12'b10111111110 		: log = 32'b00000000000000000101000101101110;
			12'b10111111111 		: log = 32'b00000000000000000101000101111010;
			12'b11000000000 		: log = 32'b00000000000000000101000110000110;
			12'b11000000001 		: log = 32'b00000000000000000101000110010001;
			12'b11000000010 		: log = 32'b00000000000000000101000110011101;
			12'b11000000011 		: log = 32'b00000000000000000101000110101001;
			12'b11000000100 		: log = 32'b00000000000000000101000110110100;
			12'b11000000101 		: log = 32'b00000000000000000101000111000000;
			12'b11000000110 		: log = 32'b00000000000000000101000111001011;
			12'b11000000111 		: log = 32'b00000000000000000101000111010111;
			12'b11000001000 		: log = 32'b00000000000000000101000111100011;
			12'b11000001001 		: log = 32'b00000000000000000101000111101110;
			12'b11000001010 		: log = 32'b00000000000000000101000111111010;
			12'b11000001011 		: log = 32'b00000000000000000101001000000110;
			12'b11000001100 		: log = 32'b00000000000000000101001000010001;
			12'b11000001101 		: log = 32'b00000000000000000101001000011101;
			12'b11000001110 		: log = 32'b00000000000000000101001000101000;
			12'b11000001111 		: log = 32'b00000000000000000101001000110100;
			12'b11000010000 		: log = 32'b00000000000000000101001001000000;
			12'b11000010001 		: log = 32'b00000000000000000101001001001011;
			12'b11000010010 		: log = 32'b00000000000000000101001001010111;
			12'b11000010011 		: log = 32'b00000000000000000101001001100010;
			12'b11000010100 		: log = 32'b00000000000000000101001001101110;
			12'b11000010101 		: log = 32'b00000000000000000101001001111010;
			12'b11000010110 		: log = 32'b00000000000000000101001010000101;
			12'b11000010111 		: log = 32'b00000000000000000101001010010001;
			12'b11000011000 		: log = 32'b00000000000000000101001010011100;
			12'b11000011001 		: log = 32'b00000000000000000101001010101000;
			12'b11000011010 		: log = 32'b00000000000000000101001010110100;
			12'b11000011011 		: log = 32'b00000000000000000101001010111111;
			12'b11000011100 		: log = 32'b00000000000000000101001011001011;
			12'b11000011101 		: log = 32'b00000000000000000101001011010110;
			12'b11000011110 		: log = 32'b00000000000000000101001011100010;
			12'b11000011111 		: log = 32'b00000000000000000101001011101101;
			12'b11000100000 		: log = 32'b00000000000000000101001011111001;
			12'b11000100001 		: log = 32'b00000000000000000101001100000101;
			12'b11000100010 		: log = 32'b00000000000000000101001100010000;
			12'b11000100011 		: log = 32'b00000000000000000101001100011100;
			12'b11000100100 		: log = 32'b00000000000000000101001100100111;
			12'b11000100101 		: log = 32'b00000000000000000101001100110011;
			12'b11000100110 		: log = 32'b00000000000000000101001100111110;
			12'b11000100111 		: log = 32'b00000000000000000101001101001010;
			12'b11000101000 		: log = 32'b00000000000000000101001101010101;
			12'b11000101001 		: log = 32'b00000000000000000101001101100001;
			12'b11000101010 		: log = 32'b00000000000000000101001101101101;
			12'b11000101011 		: log = 32'b00000000000000000101001101111000;
			12'b11000101100 		: log = 32'b00000000000000000101001110000100;
			12'b11000101101 		: log = 32'b00000000000000000101001110001111;
			12'b11000101110 		: log = 32'b00000000000000000101001110011011;
			12'b11000101111 		: log = 32'b00000000000000000101001110100110;
			12'b11000110000 		: log = 32'b00000000000000000101001110110010;
			12'b11000110001 		: log = 32'b00000000000000000101001110111101;
			12'b11000110010 		: log = 32'b00000000000000000101001111001001;
			12'b11000110011 		: log = 32'b00000000000000000101001111010100;
			12'b11000110100 		: log = 32'b00000000000000000101001111100000;
			12'b11000110101 		: log = 32'b00000000000000000101001111101100;
			12'b11000110110 		: log = 32'b00000000000000000101001111110111;
			12'b11000110111 		: log = 32'b00000000000000000101010000000011;
			12'b11000111000 		: log = 32'b00000000000000000101010000001110;
			12'b11000111001 		: log = 32'b00000000000000000101010000011010;
			12'b11000111010 		: log = 32'b00000000000000000101010000100101;
			12'b11000111011 		: log = 32'b00000000000000000101010000110001;
			12'b11000111100 		: log = 32'b00000000000000000101010000111100;
			12'b11000111101 		: log = 32'b00000000000000000101010001001000;
			12'b11000111110 		: log = 32'b00000000000000000101010001010011;
			12'b11000111111 		: log = 32'b00000000000000000101010001011111;
			12'b11001000000 		: log = 32'b00000000000000000101010001101010;
			12'b11001000001 		: log = 32'b00000000000000000101010001110110;
			12'b11001000010 		: log = 32'b00000000000000000101010010000001;
			12'b11001000011 		: log = 32'b00000000000000000101010010001101;
			12'b11001000100 		: log = 32'b00000000000000000101010010011000;
			12'b11001000101 		: log = 32'b00000000000000000101010010100100;
			12'b11001000110 		: log = 32'b00000000000000000101010010101111;
			12'b11001000111 		: log = 32'b00000000000000000101010010111011;
			12'b11001001000 		: log = 32'b00000000000000000101010011000110;
			12'b11001001001 		: log = 32'b00000000000000000101010011010010;
			12'b11001001010 		: log = 32'b00000000000000000101010011011101;
			12'b11001001011 		: log = 32'b00000000000000000101010011101001;
			12'b11001001100 		: log = 32'b00000000000000000101010011110100;
			12'b11001001101 		: log = 32'b00000000000000000101010100000000;
			12'b11001001110 		: log = 32'b00000000000000000101010100001011;
			12'b11001001111 		: log = 32'b00000000000000000101010100010111;
			12'b11001010000 		: log = 32'b00000000000000000101010100100010;
			12'b11001010001 		: log = 32'b00000000000000000101010100101110;
			12'b11001010010 		: log = 32'b00000000000000000101010100111001;
			12'b11001010011 		: log = 32'b00000000000000000101010101000100;
			12'b11001010100 		: log = 32'b00000000000000000101010101010000;
			12'b11001010101 		: log = 32'b00000000000000000101010101011011;
			12'b11001010110 		: log = 32'b00000000000000000101010101100111;
			12'b11001010111 		: log = 32'b00000000000000000101010101110010;
			12'b11001011000 		: log = 32'b00000000000000000101010101111110;
			12'b11001011001 		: log = 32'b00000000000000000101010110001001;
			12'b11001011010 		: log = 32'b00000000000000000101010110010101;
			12'b11001011011 		: log = 32'b00000000000000000101010110100000;
			12'b11001011100 		: log = 32'b00000000000000000101010110101100;
			12'b11001011101 		: log = 32'b00000000000000000101010110110111;
			12'b11001011110 		: log = 32'b00000000000000000101010111000010;
			12'b11001011111 		: log = 32'b00000000000000000101010111001110;
			12'b11001100000 		: log = 32'b00000000000000000101010111011001;
			12'b11001100001 		: log = 32'b00000000000000000101010111100101;
			12'b11001100010 		: log = 32'b00000000000000000101010111110000;
			12'b11001100011 		: log = 32'b00000000000000000101010111111100;
			12'b11001100100 		: log = 32'b00000000000000000101011000000111;
			12'b11001100101 		: log = 32'b00000000000000000101011000010011;
			12'b11001100110 		: log = 32'b00000000000000000101011000011110;
			12'b11001100111 		: log = 32'b00000000000000000101011000101001;
			12'b11001101000 		: log = 32'b00000000000000000101011000110101;
			12'b11001101001 		: log = 32'b00000000000000000101011001000000;
			12'b11001101010 		: log = 32'b00000000000000000101011001001100;
			12'b11001101011 		: log = 32'b00000000000000000101011001010111;
			12'b11001101100 		: log = 32'b00000000000000000101011001100011;
			12'b11001101101 		: log = 32'b00000000000000000101011001101110;
			12'b11001101110 		: log = 32'b00000000000000000101011001111001;
			12'b11001101111 		: log = 32'b00000000000000000101011010000101;
			12'b11001110000 		: log = 32'b00000000000000000101011010010000;
			12'b11001110001 		: log = 32'b00000000000000000101011010011100;
			12'b11001110010 		: log = 32'b00000000000000000101011010100111;
			12'b11001110011 		: log = 32'b00000000000000000101011010110010;
			12'b11001110100 		: log = 32'b00000000000000000101011010111110;
			12'b11001110101 		: log = 32'b00000000000000000101011011001001;
			12'b11001110110 		: log = 32'b00000000000000000101011011010101;
			12'b11001110111 		: log = 32'b00000000000000000101011011100000;
			12'b11001111000 		: log = 32'b00000000000000000101011011101011;
			12'b11001111001 		: log = 32'b00000000000000000101011011110111;
			12'b11001111010 		: log = 32'b00000000000000000101011100000010;
			12'b11001111011 		: log = 32'b00000000000000000101011100001110;
			12'b11001111100 		: log = 32'b00000000000000000101011100011001;
			12'b11001111101 		: log = 32'b00000000000000000101011100100100;
			12'b11001111110 		: log = 32'b00000000000000000101011100110000;
			12'b11001111111 		: log = 32'b00000000000000000101011100111011;
			12'b11010000000 		: log = 32'b00000000000000000101011101000110;
			12'b11010000001 		: log = 32'b00000000000000000101011101010010;
			12'b11010000010 		: log = 32'b00000000000000000101011101011101;
			12'b11010000011 		: log = 32'b00000000000000000101011101101001;
			12'b11010000100 		: log = 32'b00000000000000000101011101110100;
			12'b11010000101 		: log = 32'b00000000000000000101011101111111;
			12'b11010000110 		: log = 32'b00000000000000000101011110001011;
			12'b11010000111 		: log = 32'b00000000000000000101011110010110;
			12'b11010001000 		: log = 32'b00000000000000000101011110100001;
			12'b11010001001 		: log = 32'b00000000000000000101011110101101;
			12'b11010001010 		: log = 32'b00000000000000000101011110111000;
			12'b11010001011 		: log = 32'b00000000000000000101011111000100;
			12'b11010001100 		: log = 32'b00000000000000000101011111001111;
			12'b11010001101 		: log = 32'b00000000000000000101011111011010;
			12'b11010001110 		: log = 32'b00000000000000000101011111100110;
			12'b11010001111 		: log = 32'b00000000000000000101011111110001;
			12'b11010010000 		: log = 32'b00000000000000000101011111111100;
			12'b11010010001 		: log = 32'b00000000000000000101100000001000;
			12'b11010010010 		: log = 32'b00000000000000000101100000010011;
			12'b11010010011 		: log = 32'b00000000000000000101100000011110;
			12'b11010010100 		: log = 32'b00000000000000000101100000101010;
			12'b11010010101 		: log = 32'b00000000000000000101100000110101;
			12'b11010010110 		: log = 32'b00000000000000000101100001000000;
			12'b11010010111 		: log = 32'b00000000000000000101100001001100;
			12'b11010011000 		: log = 32'b00000000000000000101100001010111;
			12'b11010011001 		: log = 32'b00000000000000000101100001100010;
			12'b11010011010 		: log = 32'b00000000000000000101100001101110;
			12'b11010011011 		: log = 32'b00000000000000000101100001111001;
			12'b11010011100 		: log = 32'b00000000000000000101100010000100;
			12'b11010011101 		: log = 32'b00000000000000000101100010010000;
			12'b11010011110 		: log = 32'b00000000000000000101100010011011;
			12'b11010011111 		: log = 32'b00000000000000000101100010100110;
			12'b11010100000 		: log = 32'b00000000000000000101100010110010;
			12'b11010100001 		: log = 32'b00000000000000000101100010111101;
			12'b11010100010 		: log = 32'b00000000000000000101100011001000;
			12'b11010100011 		: log = 32'b00000000000000000101100011010011;
			12'b11010100100 		: log = 32'b00000000000000000101100011011111;
			12'b11010100101 		: log = 32'b00000000000000000101100011101010;
			12'b11010100110 		: log = 32'b00000000000000000101100011110101;
			12'b11010100111 		: log = 32'b00000000000000000101100100000001;
			12'b11010101000 		: log = 32'b00000000000000000101100100001100;
			12'b11010101001 		: log = 32'b00000000000000000101100100010111;
			12'b11010101010 		: log = 32'b00000000000000000101100100100011;
			12'b11010101011 		: log = 32'b00000000000000000101100100101110;
			12'b11010101100 		: log = 32'b00000000000000000101100100111001;
			12'b11010101101 		: log = 32'b00000000000000000101100101000100;
			12'b11010101110 		: log = 32'b00000000000000000101100101010000;
			12'b11010101111 		: log = 32'b00000000000000000101100101011011;
			12'b11010110000 		: log = 32'b00000000000000000101100101100110;
			12'b11010110001 		: log = 32'b00000000000000000101100101110010;
			12'b11010110010 		: log = 32'b00000000000000000101100101111101;
			12'b11010110011 		: log = 32'b00000000000000000101100110001000;
			12'b11010110100 		: log = 32'b00000000000000000101100110010011;
			12'b11010110101 		: log = 32'b00000000000000000101100110011111;
			12'b11010110110 		: log = 32'b00000000000000000101100110101010;
			12'b11010110111 		: log = 32'b00000000000000000101100110110101;
			12'b11010111000 		: log = 32'b00000000000000000101100111000001;
			12'b11010111001 		: log = 32'b00000000000000000101100111001100;
			12'b11010111010 		: log = 32'b00000000000000000101100111010111;
			12'b11010111011 		: log = 32'b00000000000000000101100111100010;
			12'b11010111100 		: log = 32'b00000000000000000101100111101110;
			12'b11010111101 		: log = 32'b00000000000000000101100111111001;
			12'b11010111110 		: log = 32'b00000000000000000101101000000100;
			12'b11010111111 		: log = 32'b00000000000000000101101000001111;
			12'b11011000000 		: log = 32'b00000000000000000101101000011011;
			12'b11011000001 		: log = 32'b00000000000000000101101000100110;
			12'b11011000010 		: log = 32'b00000000000000000101101000110001;
			12'b11011000011 		: log = 32'b00000000000000000101101000111100;
			12'b11011000100 		: log = 32'b00000000000000000101101001001000;
			12'b11011000101 		: log = 32'b00000000000000000101101001010011;
			12'b11011000110 		: log = 32'b00000000000000000101101001011110;
			12'b11011000111 		: log = 32'b00000000000000000101101001101001;
			12'b11011001000 		: log = 32'b00000000000000000101101001110101;
			12'b11011001001 		: log = 32'b00000000000000000101101010000000;
			12'b11011001010 		: log = 32'b00000000000000000101101010001011;
			12'b11011001011 		: log = 32'b00000000000000000101101010010110;
			12'b11011001100 		: log = 32'b00000000000000000101101010100010;
			12'b11011001101 		: log = 32'b00000000000000000101101010101101;
			12'b11011001110 		: log = 32'b00000000000000000101101010111000;
			12'b11011001111 		: log = 32'b00000000000000000101101011000011;
			12'b11011010000 		: log = 32'b00000000000000000101101011001110;
			12'b11011010001 		: log = 32'b00000000000000000101101011011010;
			12'b11011010010 		: log = 32'b00000000000000000101101011100101;
			12'b11011010011 		: log = 32'b00000000000000000101101011110000;
			12'b11011010100 		: log = 32'b00000000000000000101101011111011;
			12'b11011010101 		: log = 32'b00000000000000000101101100000111;
			12'b11011010110 		: log = 32'b00000000000000000101101100010010;
			12'b11011010111 		: log = 32'b00000000000000000101101100011101;
			12'b11011011000 		: log = 32'b00000000000000000101101100101000;
			12'b11011011001 		: log = 32'b00000000000000000101101100110011;
			12'b11011011010 		: log = 32'b00000000000000000101101100111111;
			12'b11011011011 		: log = 32'b00000000000000000101101101001010;
			12'b11011011100 		: log = 32'b00000000000000000101101101010101;
			12'b11011011101 		: log = 32'b00000000000000000101101101100000;
			12'b11011011110 		: log = 32'b00000000000000000101101101101011;
			12'b11011011111 		: log = 32'b00000000000000000101101101110111;
			12'b11011100000 		: log = 32'b00000000000000000101101110000010;
			12'b11011100001 		: log = 32'b00000000000000000101101110001101;
			12'b11011100010 		: log = 32'b00000000000000000101101110011000;
			12'b11011100011 		: log = 32'b00000000000000000101101110100011;
			12'b11011100100 		: log = 32'b00000000000000000101101110101110;
			12'b11011100101 		: log = 32'b00000000000000000101101110111010;
			12'b11011100110 		: log = 32'b00000000000000000101101111000101;
			12'b11011100111 		: log = 32'b00000000000000000101101111010000;
			12'b11011101000 		: log = 32'b00000000000000000101101111011011;
			12'b11011101001 		: log = 32'b00000000000000000101101111100110;
			12'b11011101010 		: log = 32'b00000000000000000101101111110010;
			12'b11011101011 		: log = 32'b00000000000000000101101111111101;
			12'b11011101100 		: log = 32'b00000000000000000101110000001000;
			12'b11011101101 		: log = 32'b00000000000000000101110000010011;
			12'b11011101110 		: log = 32'b00000000000000000101110000011110;
			12'b11011101111 		: log = 32'b00000000000000000101110000101001;
			12'b11011110000 		: log = 32'b00000000000000000101110000110101;
			12'b11011110001 		: log = 32'b00000000000000000101110001000000;
			12'b11011110010 		: log = 32'b00000000000000000101110001001011;
			12'b11011110011 		: log = 32'b00000000000000000101110001010110;
			12'b11011110100 		: log = 32'b00000000000000000101110001100001;
			12'b11011110101 		: log = 32'b00000000000000000101110001101100;
			12'b11011110110 		: log = 32'b00000000000000000101110001110111;
			12'b11011110111 		: log = 32'b00000000000000000101110010000011;
			12'b11011111000 		: log = 32'b00000000000000000101110010001110;
			12'b11011111001 		: log = 32'b00000000000000000101110010011001;
			12'b11011111010 		: log = 32'b00000000000000000101110010100100;
			12'b11011111011 		: log = 32'b00000000000000000101110010101111;
			12'b11011111100 		: log = 32'b00000000000000000101110010111010;
			12'b11011111101 		: log = 32'b00000000000000000101110011000101;
			12'b11011111110 		: log = 32'b00000000000000000101110011010001;
			12'b11011111111 		: log = 32'b00000000000000000101110011011100;
			12'b11100000000 		: log = 32'b00000000000000000101110011100111;
			12'b11100000001 		: log = 32'b00000000000000000101110011110010;
			12'b11100000010 		: log = 32'b00000000000000000101110011111101;
			12'b11100000011 		: log = 32'b00000000000000000101110100001000;
			12'b11100000100 		: log = 32'b00000000000000000101110100010011;
			12'b11100000101 		: log = 32'b00000000000000000101110100011111;
			12'b11100000110 		: log = 32'b00000000000000000101110100101010;
			12'b11100000111 		: log = 32'b00000000000000000101110100110101;
			12'b11100001000 		: log = 32'b00000000000000000101110101000000;
			12'b11100001001 		: log = 32'b00000000000000000101110101001011;
			12'b11100001010 		: log = 32'b00000000000000000101110101010110;
			12'b11100001011 		: log = 32'b00000000000000000101110101100001;
			12'b11100001100 		: log = 32'b00000000000000000101110101101100;
			12'b11100001101 		: log = 32'b00000000000000000101110101110111;
			12'b11100001110 		: log = 32'b00000000000000000101110110000011;
			12'b11100001111 		: log = 32'b00000000000000000101110110001110;
			12'b11100010000 		: log = 32'b00000000000000000101110110011001;
			12'b11100010001 		: log = 32'b00000000000000000101110110100100;
			12'b11100010010 		: log = 32'b00000000000000000101110110101111;
			12'b11100010011 		: log = 32'b00000000000000000101110110111010;
			12'b11100010100 		: log = 32'b00000000000000000101110111000101;
			12'b11100010101 		: log = 32'b00000000000000000101110111010000;
			12'b11100010110 		: log = 32'b00000000000000000101110111011011;
			12'b11100010111 		: log = 32'b00000000000000000101110111100110;
			12'b11100011000 		: log = 32'b00000000000000000101110111110001;
			12'b11100011001 		: log = 32'b00000000000000000101110111111101;
			12'b11100011010 		: log = 32'b00000000000000000101111000001000;
			12'b11100011011 		: log = 32'b00000000000000000101111000010011;
			12'b11100011100 		: log = 32'b00000000000000000101111000011110;
			12'b11100011101 		: log = 32'b00000000000000000101111000101001;
			12'b11100011110 		: log = 32'b00000000000000000101111000110100;
			12'b11100011111 		: log = 32'b00000000000000000101111000111111;
			12'b11100100000 		: log = 32'b00000000000000000101111001001010;
			12'b11100100001 		: log = 32'b00000000000000000101111001010101;
			12'b11100100010 		: log = 32'b00000000000000000101111001100000;
			12'b11100100011 		: log = 32'b00000000000000000101111001101011;
			12'b11100100100 		: log = 32'b00000000000000000101111001110110;
			12'b11100100101 		: log = 32'b00000000000000000101111010000001;
			12'b11100100110 		: log = 32'b00000000000000000101111010001100;
			12'b11100100111 		: log = 32'b00000000000000000101111010011000;
			12'b11100101000 		: log = 32'b00000000000000000101111010100011;
			12'b11100101001 		: log = 32'b00000000000000000101111010101110;
			12'b11100101010 		: log = 32'b00000000000000000101111010111001;
			12'b11100101011 		: log = 32'b00000000000000000101111011000100;
			12'b11100101100 		: log = 32'b00000000000000000101111011001111;
			12'b11100101101 		: log = 32'b00000000000000000101111011011010;
			12'b11100101110 		: log = 32'b00000000000000000101111011100101;
			12'b11100101111 		: log = 32'b00000000000000000101111011110000;
			12'b11100110000 		: log = 32'b00000000000000000101111011111011;
			12'b11100110001 		: log = 32'b00000000000000000101111100000110;
			12'b11100110010 		: log = 32'b00000000000000000101111100010001;
			12'b11100110011 		: log = 32'b00000000000000000101111100011100;
			12'b11100110100 		: log = 32'b00000000000000000101111100100111;
			12'b11100110101 		: log = 32'b00000000000000000101111100110010;
			12'b11100110110 		: log = 32'b00000000000000000101111100111101;
			12'b11100110111 		: log = 32'b00000000000000000101111101001000;
			12'b11100111000 		: log = 32'b00000000000000000101111101010011;
			12'b11100111001 		: log = 32'b00000000000000000101111101011110;
			12'b11100111010 		: log = 32'b00000000000000000101111101101001;
			12'b11100111011 		: log = 32'b00000000000000000101111101110100;
			12'b11100111100 		: log = 32'b00000000000000000101111101111111;
			12'b11100111101 		: log = 32'b00000000000000000101111110001010;
			12'b11100111110 		: log = 32'b00000000000000000101111110010101;
			12'b11100111111 		: log = 32'b00000000000000000101111110100000;
			12'b11101000000 		: log = 32'b00000000000000000101111110101011;
			12'b11101000001 		: log = 32'b00000000000000000101111110110110;
			12'b11101000010 		: log = 32'b00000000000000000101111111000001;
			12'b11101000011 		: log = 32'b00000000000000000101111111001100;
			12'b11101000100 		: log = 32'b00000000000000000101111111010111;
			12'b11101000101 		: log = 32'b00000000000000000101111111100010;
			12'b11101000110 		: log = 32'b00000000000000000101111111101101;
			12'b11101000111 		: log = 32'b00000000000000000101111111111000;
			12'b11101001000 		: log = 32'b00000000000000000110000000000011;
			12'b11101001001 		: log = 32'b00000000000000000110000000001110;
			12'b11101001010 		: log = 32'b00000000000000000110000000011001;
			12'b11101001011 		: log = 32'b00000000000000000110000000100100;
			12'b11101001100 		: log = 32'b00000000000000000110000000101111;
			12'b11101001101 		: log = 32'b00000000000000000110000000111010;
			12'b11101001110 		: log = 32'b00000000000000000110000001000101;
			12'b11101001111 		: log = 32'b00000000000000000110000001010000;
			12'b11101010000 		: log = 32'b00000000000000000110000001011011;
			12'b11101010001 		: log = 32'b00000000000000000110000001100110;
			12'b11101010010 		: log = 32'b00000000000000000110000001110001;
			12'b11101010011 		: log = 32'b00000000000000000110000001111100;
			12'b11101010100 		: log = 32'b00000000000000000110000010000111;
			12'b11101010101 		: log = 32'b00000000000000000110000010010010;
			12'b11101010110 		: log = 32'b00000000000000000110000010011101;
			12'b11101010111 		: log = 32'b00000000000000000110000010101000;
			12'b11101011000 		: log = 32'b00000000000000000110000010110011;
			12'b11101011001 		: log = 32'b00000000000000000110000010111110;
			12'b11101011010 		: log = 32'b00000000000000000110000011001001;
			12'b11101011011 		: log = 32'b00000000000000000110000011010100;
			12'b11101011100 		: log = 32'b00000000000000000110000011011111;
			12'b11101011101 		: log = 32'b00000000000000000110000011101010;
			12'b11101011110 		: log = 32'b00000000000000000110000011110101;
			12'b11101011111 		: log = 32'b00000000000000000110000100000000;
			12'b11101100000 		: log = 32'b00000000000000000110000100001011;
			12'b11101100001 		: log = 32'b00000000000000000110000100010110;
			12'b11101100010 		: log = 32'b00000000000000000110000100100001;
			12'b11101100011 		: log = 32'b00000000000000000110000100101100;
			12'b11101100100 		: log = 32'b00000000000000000110000100110111;
			12'b11101100101 		: log = 32'b00000000000000000110000101000010;
			12'b11101100110 		: log = 32'b00000000000000000110000101001100;
			12'b11101100111 		: log = 32'b00000000000000000110000101010111;
			12'b11101101000 		: log = 32'b00000000000000000110000101100010;
			12'b11101101001 		: log = 32'b00000000000000000110000101101101;
			12'b11101101010 		: log = 32'b00000000000000000110000101111000;
			12'b11101101011 		: log = 32'b00000000000000000110000110000011;
			12'b11101101100 		: log = 32'b00000000000000000110000110001110;
			12'b11101101101 		: log = 32'b00000000000000000110000110011001;
			12'b11101101110 		: log = 32'b00000000000000000110000110100100;
			12'b11101101111 		: log = 32'b00000000000000000110000110101111;
			12'b11101110000 		: log = 32'b00000000000000000110000110111010;
			12'b11101110001 		: log = 32'b00000000000000000110000111000101;
			12'b11101110010 		: log = 32'b00000000000000000110000111010000;
			12'b11101110011 		: log = 32'b00000000000000000110000111011011;
			12'b11101110100 		: log = 32'b00000000000000000110000111100101;
			12'b11101110101 		: log = 32'b00000000000000000110000111110000;
			12'b11101110110 		: log = 32'b00000000000000000110000111111011;
			12'b11101110111 		: log = 32'b00000000000000000110001000000110;
			12'b11101111000 		: log = 32'b00000000000000000110001000010001;
			12'b11101111001 		: log = 32'b00000000000000000110001000011100;
			12'b11101111010 		: log = 32'b00000000000000000110001000100111;
			12'b11101111011 		: log = 32'b00000000000000000110001000110010;
			12'b11101111100 		: log = 32'b00000000000000000110001000111101;
			12'b11101111101 		: log = 32'b00000000000000000110001001001000;
			12'b11101111110 		: log = 32'b00000000000000000110001001010011;
			12'b11101111111 		: log = 32'b00000000000000000110001001011101;
			12'b11110000000 		: log = 32'b00000000000000000110001001101000;
			12'b11110000001 		: log = 32'b00000000000000000110001001110011;
			12'b11110000010 		: log = 32'b00000000000000000110001001111110;
			12'b11110000011 		: log = 32'b00000000000000000110001010001001;
			12'b11110000100 		: log = 32'b00000000000000000110001010010100;
			12'b11110000101 		: log = 32'b00000000000000000110001010011111;
			12'b11110000110 		: log = 32'b00000000000000000110001010101010;
			12'b11110000111 		: log = 32'b00000000000000000110001010110101;
			12'b11110001000 		: log = 32'b00000000000000000110001010111111;
			12'b11110001001 		: log = 32'b00000000000000000110001011001010;
			12'b11110001010 		: log = 32'b00000000000000000110001011010101;
			12'b11110001011 		: log = 32'b00000000000000000110001011100000;
			12'b11110001100 		: log = 32'b00000000000000000110001011101011;
			12'b11110001101 		: log = 32'b00000000000000000110001011110110;
			12'b11110001110 		: log = 32'b00000000000000000110001100000001;
			12'b11110001111 		: log = 32'b00000000000000000110001100001100;
			12'b11110010000 		: log = 32'b00000000000000000110001100010110;
			12'b11110010001 		: log = 32'b00000000000000000110001100100001;
			12'b11110010010 		: log = 32'b00000000000000000110001100101100;
			12'b11110010011 		: log = 32'b00000000000000000110001100110111;
			12'b11110010100 		: log = 32'b00000000000000000110001101000010;
			12'b11110010101 		: log = 32'b00000000000000000110001101001101;
			12'b11110010110 		: log = 32'b00000000000000000110001101011000;
			12'b11110010111 		: log = 32'b00000000000000000110001101100010;
			12'b11110011000 		: log = 32'b00000000000000000110001101101101;
			12'b11110011001 		: log = 32'b00000000000000000110001101111000;
			12'b11110011010 		: log = 32'b00000000000000000110001110000011;
			12'b11110011011 		: log = 32'b00000000000000000110001110001110;
			12'b11110011100 		: log = 32'b00000000000000000110001110011001;
			12'b11110011101 		: log = 32'b00000000000000000110001110100011;
			12'b11110011110 		: log = 32'b00000000000000000110001110101110;
			12'b11110011111 		: log = 32'b00000000000000000110001110111001;
			12'b11110100000 		: log = 32'b00000000000000000110001111000100;
			12'b11110100001 		: log = 32'b00000000000000000110001111001111;
			12'b11110100010 		: log = 32'b00000000000000000110001111011010;
			12'b11110100011 		: log = 32'b00000000000000000110001111100100;
			12'b11110100100 		: log = 32'b00000000000000000110001111101111;
			12'b11110100101 		: log = 32'b00000000000000000110001111111010;
			12'b11110100110 		: log = 32'b00000000000000000110010000000101;
			12'b11110100111 		: log = 32'b00000000000000000110010000010000;
			12'b11110101000 		: log = 32'b00000000000000000110010000011011;
			12'b11110101001 		: log = 32'b00000000000000000110010000100101;
			12'b11110101010 		: log = 32'b00000000000000000110010000110000;
			12'b11110101011 		: log = 32'b00000000000000000110010000111011;
			12'b11110101100 		: log = 32'b00000000000000000110010001000110;
			12'b11110101101 		: log = 32'b00000000000000000110010001010001;
			12'b11110101110 		: log = 32'b00000000000000000110010001011100;
			12'b11110101111 		: log = 32'b00000000000000000110010001100110;
			12'b11110110000 		: log = 32'b00000000000000000110010001110001;
			12'b11110110001 		: log = 32'b00000000000000000110010001111100;
			12'b11110110010 		: log = 32'b00000000000000000110010010000111;
			12'b11110110011 		: log = 32'b00000000000000000110010010010010;
			12'b11110110100 		: log = 32'b00000000000000000110010010011100;
			12'b11110110101 		: log = 32'b00000000000000000110010010100111;
			12'b11110110110 		: log = 32'b00000000000000000110010010110010;
			12'b11110110111 		: log = 32'b00000000000000000110010010111101;
			12'b11110111000 		: log = 32'b00000000000000000110010011001000;
			12'b11110111001 		: log = 32'b00000000000000000110010011010010;
			12'b11110111010 		: log = 32'b00000000000000000110010011011101;
			12'b11110111011 		: log = 32'b00000000000000000110010011101000;
			12'b11110111100 		: log = 32'b00000000000000000110010011110011;
			12'b11110111101 		: log = 32'b00000000000000000110010011111101;
			12'b11110111110 		: log = 32'b00000000000000000110010100001000;
			12'b11110111111 		: log = 32'b00000000000000000110010100010011;
			12'b11111000000 		: log = 32'b00000000000000000110010100011110;
			12'b11111000001 		: log = 32'b00000000000000000110010100101001;
			12'b11111000010 		: log = 32'b00000000000000000110010100110011;
			12'b11111000011 		: log = 32'b00000000000000000110010100111110;
			12'b11111000100 		: log = 32'b00000000000000000110010101001001;
			12'b11111000101 		: log = 32'b00000000000000000110010101010100;
			12'b11111000110 		: log = 32'b00000000000000000110010101011110;
			12'b11111000111 		: log = 32'b00000000000000000110010101101001;
			12'b11111001000 		: log = 32'b00000000000000000110010101110100;
			12'b11111001001 		: log = 32'b00000000000000000110010101111111;
			12'b11111001010 		: log = 32'b00000000000000000110010110001010;
			12'b11111001011 		: log = 32'b00000000000000000110010110010100;
			12'b11111001100 		: log = 32'b00000000000000000110010110011111;
			12'b11111001101 		: log = 32'b00000000000000000110010110101010;
			12'b11111001110 		: log = 32'b00000000000000000110010110110101;
			12'b11111001111 		: log = 32'b00000000000000000110010110111111;
			12'b11111010000 		: log = 32'b00000000000000000110010111001010;
			12'b11111010001 		: log = 32'b00000000000000000110010111010101;
			12'b11111010010 		: log = 32'b00000000000000000110010111100000;
			12'b11111010011 		: log = 32'b00000000000000000110010111101010;
			12'b11111010100 		: log = 32'b00000000000000000110010111110101;
			12'b11111010101 		: log = 32'b00000000000000000110011000000000;
			12'b11111010110 		: log = 32'b00000000000000000110011000001011;
			12'b11111010111 		: log = 32'b00000000000000000110011000010101;
			12'b11111011000 		: log = 32'b00000000000000000110011000100000;
			12'b11111011001 		: log = 32'b00000000000000000110011000101011;
			12'b11111011010 		: log = 32'b00000000000000000110011000110101;
			12'b11111011011 		: log = 32'b00000000000000000110011001000000;
			12'b11111011100 		: log = 32'b00000000000000000110011001001011;
			12'b11111011101 		: log = 32'b00000000000000000110011001010110;
			12'b11111011110 		: log = 32'b00000000000000000110011001100000;
			12'b11111011111 		: log = 32'b00000000000000000110011001101011;
			12'b11111100000 		: log = 32'b00000000000000000110011001110110;
			12'b11111100001 		: log = 32'b00000000000000000110011010000001;
			12'b11111100010 		: log = 32'b00000000000000000110011010001011;
			12'b11111100011 		: log = 32'b00000000000000000110011010010110;
			12'b11111100100 		: log = 32'b00000000000000000110011010100001;
			12'b11111100101 		: log = 32'b00000000000000000110011010101011;
			12'b11111100110 		: log = 32'b00000000000000000110011010110110;
			12'b11111100111 		: log = 32'b00000000000000000110011011000001;
			12'b11111101000 		: log = 32'b00000000000000000110011011001100;
			12'b11111101001 		: log = 32'b00000000000000000110011011010110;
			12'b11111101010 		: log = 32'b00000000000000000110011011100001;
			12'b11111101011 		: log = 32'b00000000000000000110011011101100;
			12'b11111101100 		: log = 32'b00000000000000000110011011110110;
			12'b11111101101 		: log = 32'b00000000000000000110011100000001;
			12'b11111101110 		: log = 32'b00000000000000000110011100001100;
			12'b11111101111 		: log = 32'b00000000000000000110011100010110;
			12'b11111110000 		: log = 32'b00000000000000000110011100100001;
			12'b11111110001 		: log = 32'b00000000000000000110011100101100;
			12'b11111110010 		: log = 32'b00000000000000000110011100110111;
			12'b11111110011 		: log = 32'b00000000000000000110011101000001;
			12'b11111110100 		: log = 32'b00000000000000000110011101001100;
			12'b11111110101 		: log = 32'b00000000000000000110011101010111;
			12'b11111110110 		: log = 32'b00000000000000000110011101100001;
			12'b11111110111 		: log = 32'b00000000000000000110011101101100;
			12'b11111111000 		: log = 32'b00000000000000000110011101110111;
			12'b11111111001 		: log = 32'b00000000000000000110011110000001;
			12'b11111111010 		: log = 32'b00000000000000000110011110001100;
			12'b11111111011 		: log = 32'b00000000000000000110011110010111;
			12'b11111111100 		: log = 32'b00000000000000000110011110100001;
			12'b11111111101 		: log = 32'b00000000000000000110011110101100;
			12'b11111111110 		: log = 32'b00000000000000000110011110110111;
			12'b11111111111 		: log = 32'b00000000000000000110011111000001;
			12'b100000000000 		: log = 32'b00000000000000000110011111001100;
			12'b100000000001 		: log = 32'b00000000000000000110011111010111;
			12'b100000000010 		: log = 32'b00000000000000000110011111100001;
			12'b100000000011 		: log = 32'b00000000000000000110011111101100;
			12'b100000000100 		: log = 32'b00000000000000000110011111110111;
			12'b100000000101 		: log = 32'b00000000000000000110100000000001;
			12'b100000000110 		: log = 32'b00000000000000000110100000001100;
			12'b100000000111 		: log = 32'b00000000000000000110100000010111;
			12'b100000001000 		: log = 32'b00000000000000000110100000100001;
			12'b100000001001 		: log = 32'b00000000000000000110100000101100;
			12'b100000001010 		: log = 32'b00000000000000000110100000110111;
			12'b100000001011 		: log = 32'b00000000000000000110100001000001;
			12'b100000001100 		: log = 32'b00000000000000000110100001001100;
			12'b100000001101 		: log = 32'b00000000000000000110100001010111;
			12'b100000001110 		: log = 32'b00000000000000000110100001100001;
			12'b100000001111 		: log = 32'b00000000000000000110100001101100;
			12'b100000010000 		: log = 32'b00000000000000000110100001110111;
			12'b100000010001 		: log = 32'b00000000000000000110100010000001;
			12'b100000010010 		: log = 32'b00000000000000000110100010001100;
			12'b100000010011 		: log = 32'b00000000000000000110100010010110;
			12'b100000010100 		: log = 32'b00000000000000000110100010100001;
			12'b100000010101 		: log = 32'b00000000000000000110100010101100;
			12'b100000010110 		: log = 32'b00000000000000000110100010110110;
			12'b100000010111 		: log = 32'b00000000000000000110100011000001;
			12'b100000011000 		: log = 32'b00000000000000000110100011001100;
			12'b100000011001 		: log = 32'b00000000000000000110100011010110;
			12'b100000011010 		: log = 32'b00000000000000000110100011100001;
			12'b100000011011 		: log = 32'b00000000000000000110100011101011;
			12'b100000011100 		: log = 32'b00000000000000000110100011110110;
			12'b100000011101 		: log = 32'b00000000000000000110100100000001;
			12'b100000011110 		: log = 32'b00000000000000000110100100001011;
			12'b100000011111 		: log = 32'b00000000000000000110100100010110;
			12'b100000100000 		: log = 32'b00000000000000000110100100100001;
			12'b100000100001 		: log = 32'b00000000000000000110100100101011;
			12'b100000100010 		: log = 32'b00000000000000000110100100110110;
			12'b100000100011 		: log = 32'b00000000000000000110100101000000;
			12'b100000100100 		: log = 32'b00000000000000000110100101001011;
			12'b100000100101 		: log = 32'b00000000000000000110100101010110;
			12'b100000100110 		: log = 32'b00000000000000000110100101100000;
			12'b100000100111 		: log = 32'b00000000000000000110100101101011;
			12'b100000101000 		: log = 32'b00000000000000000110100101110101;
			12'b100000101001 		: log = 32'b00000000000000000110100110000000;
			12'b100000101010 		: log = 32'b00000000000000000110100110001011;
			12'b100000101011 		: log = 32'b00000000000000000110100110010101;
			12'b100000101100 		: log = 32'b00000000000000000110100110100000;
			12'b100000101101 		: log = 32'b00000000000000000110100110101010;
			12'b100000101110 		: log = 32'b00000000000000000110100110110101;
			12'b100000101111 		: log = 32'b00000000000000000110100110111111;
			12'b100000110000 		: log = 32'b00000000000000000110100111001010;
			12'b100000110001 		: log = 32'b00000000000000000110100111010101;
			12'b100000110010 		: log = 32'b00000000000000000110100111011111;
			12'b100000110011 		: log = 32'b00000000000000000110100111101010;
			12'b100000110100 		: log = 32'b00000000000000000110100111110100;
			12'b100000110101 		: log = 32'b00000000000000000110100111111111;
			12'b100000110110 		: log = 32'b00000000000000000110101000001010;
			12'b100000110111 		: log = 32'b00000000000000000110101000010100;
			12'b100000111000 		: log = 32'b00000000000000000110101000011111;
			12'b100000111001 		: log = 32'b00000000000000000110101000101001;
			12'b100000111010 		: log = 32'b00000000000000000110101000110100;
			12'b100000111011 		: log = 32'b00000000000000000110101000111110;
			12'b100000111100 		: log = 32'b00000000000000000110101001001001;
			12'b100000111101 		: log = 32'b00000000000000000110101001010100;
			12'b100000111110 		: log = 32'b00000000000000000110101001011110;
			12'b100000111111 		: log = 32'b00000000000000000110101001101001;
			12'b100001000000 		: log = 32'b00000000000000000110101001110011;
			12'b100001000001 		: log = 32'b00000000000000000110101001111110;
			12'b100001000010 		: log = 32'b00000000000000000110101010001000;
			12'b100001000011 		: log = 32'b00000000000000000110101010010011;
			12'b100001000100 		: log = 32'b00000000000000000110101010011101;
			12'b100001000101 		: log = 32'b00000000000000000110101010101000;
			12'b100001000110 		: log = 32'b00000000000000000110101010110011;
			12'b100001000111 		: log = 32'b00000000000000000110101010111101;
			12'b100001001000 		: log = 32'b00000000000000000110101011001000;
			12'b100001001001 		: log = 32'b00000000000000000110101011010010;
			12'b100001001010 		: log = 32'b00000000000000000110101011011101;
			12'b100001001011 		: log = 32'b00000000000000000110101011100111;
			12'b100001001100 		: log = 32'b00000000000000000110101011110010;
			12'b100001001101 		: log = 32'b00000000000000000110101011111100;
			12'b100001001110 		: log = 32'b00000000000000000110101100000111;
			12'b100001001111 		: log = 32'b00000000000000000110101100010001;
			12'b100001010000 		: log = 32'b00000000000000000110101100011100;
			12'b100001010001 		: log = 32'b00000000000000000110101100100110;
			12'b100001010010 		: log = 32'b00000000000000000110101100110001;
			12'b100001010011 		: log = 32'b00000000000000000110101100111011;
			12'b100001010100 		: log = 32'b00000000000000000110101101000110;
			12'b100001010101 		: log = 32'b00000000000000000110101101010001;
			12'b100001010110 		: log = 32'b00000000000000000110101101011011;
			12'b100001010111 		: log = 32'b00000000000000000110101101100110;
			12'b100001011000 		: log = 32'b00000000000000000110101101110000;
			12'b100001011001 		: log = 32'b00000000000000000110101101111011;
			12'b100001011010 		: log = 32'b00000000000000000110101110000101;
			12'b100001011011 		: log = 32'b00000000000000000110101110010000;
			12'b100001011100 		: log = 32'b00000000000000000110101110011010;
			12'b100001011101 		: log = 32'b00000000000000000110101110100101;
			12'b100001011110 		: log = 32'b00000000000000000110101110101111;
			12'b100001011111 		: log = 32'b00000000000000000110101110111010;
			12'b100001100000 		: log = 32'b00000000000000000110101111000100;
			12'b100001100001 		: log = 32'b00000000000000000110101111001111;
			12'b100001100010 		: log = 32'b00000000000000000110101111011001;
			12'b100001100011 		: log = 32'b00000000000000000110101111100100;
			12'b100001100100 		: log = 32'b00000000000000000110101111101110;
			12'b100001100101 		: log = 32'b00000000000000000110101111111001;
			12'b100001100110 		: log = 32'b00000000000000000110110000000011;
			12'b100001100111 		: log = 32'b00000000000000000110110000001110;
			12'b100001101000 		: log = 32'b00000000000000000110110000011000;
			12'b100001101001 		: log = 32'b00000000000000000110110000100011;
			12'b100001101010 		: log = 32'b00000000000000000110110000101101;
			12'b100001101011 		: log = 32'b00000000000000000110110000111000;
			12'b100001101100 		: log = 32'b00000000000000000110110001000010;
			12'b100001101101 		: log = 32'b00000000000000000110110001001101;
			12'b100001101110 		: log = 32'b00000000000000000110110001010111;
			12'b100001101111 		: log = 32'b00000000000000000110110001100001;
			12'b100001110000 		: log = 32'b00000000000000000110110001101100;
			12'b100001110001 		: log = 32'b00000000000000000110110001110110;
			12'b100001110010 		: log = 32'b00000000000000000110110010000001;
			12'b100001110011 		: log = 32'b00000000000000000110110010001011;
			12'b100001110100 		: log = 32'b00000000000000000110110010010110;
			12'b100001110101 		: log = 32'b00000000000000000110110010100000;
			12'b100001110110 		: log = 32'b00000000000000000110110010101011;
			12'b100001110111 		: log = 32'b00000000000000000110110010110101;
			12'b100001111000 		: log = 32'b00000000000000000110110011000000;
			12'b100001111001 		: log = 32'b00000000000000000110110011001010;
			12'b100001111010 		: log = 32'b00000000000000000110110011010101;
			12'b100001111011 		: log = 32'b00000000000000000110110011011111;
			12'b100001111100 		: log = 32'b00000000000000000110110011101010;
			12'b100001111101 		: log = 32'b00000000000000000110110011110100;
			12'b100001111110 		: log = 32'b00000000000000000110110011111110;
			12'b100001111111 		: log = 32'b00000000000000000110110100001001;
			12'b100010000000 		: log = 32'b00000000000000000110110100010011;
			12'b100010000001 		: log = 32'b00000000000000000110110100011110;
			12'b100010000010 		: log = 32'b00000000000000000110110100101000;
			12'b100010000011 		: log = 32'b00000000000000000110110100110011;
			12'b100010000100 		: log = 32'b00000000000000000110110100111101;
			12'b100010000101 		: log = 32'b00000000000000000110110101001000;
			12'b100010000110 		: log = 32'b00000000000000000110110101010010;
			12'b100010000111 		: log = 32'b00000000000000000110110101011100;
			12'b100010001000 		: log = 32'b00000000000000000110110101100111;
			12'b100010001001 		: log = 32'b00000000000000000110110101110001;
			12'b100010001010 		: log = 32'b00000000000000000110110101111100;
			12'b100010001011 		: log = 32'b00000000000000000110110110000110;
			12'b100010001100 		: log = 32'b00000000000000000110110110010001;
			12'b100010001101 		: log = 32'b00000000000000000110110110011011;
			12'b100010001110 		: log = 32'b00000000000000000110110110100101;
			12'b100010001111 		: log = 32'b00000000000000000110110110110000;
			12'b100010010000 		: log = 32'b00000000000000000110110110111010;
			12'b100010010001 		: log = 32'b00000000000000000110110111000101;
			12'b100010010010 		: log = 32'b00000000000000000110110111001111;
			12'b100010010011 		: log = 32'b00000000000000000110110111011010;
			12'b100010010100 		: log = 32'b00000000000000000110110111100100;
			12'b100010010101 		: log = 32'b00000000000000000110110111101110;
			12'b100010010110 		: log = 32'b00000000000000000110110111111001;
			12'b100010010111 		: log = 32'b00000000000000000110111000000011;
			12'b100010011000 		: log = 32'b00000000000000000110111000001110;
			12'b100010011001 		: log = 32'b00000000000000000110111000011000;
			12'b100010011010 		: log = 32'b00000000000000000110111000100010;
			12'b100010011011 		: log = 32'b00000000000000000110111000101101;
			12'b100010011100 		: log = 32'b00000000000000000110111000110111;
			12'b100010011101 		: log = 32'b00000000000000000110111001000010;
			12'b100010011110 		: log = 32'b00000000000000000110111001001100;
			12'b100010011111 		: log = 32'b00000000000000000110111001010110;
			12'b100010100000 		: log = 32'b00000000000000000110111001100001;
			12'b100010100001 		: log = 32'b00000000000000000110111001101011;
			12'b100010100010 		: log = 32'b00000000000000000110111001110110;
			12'b100010100011 		: log = 32'b00000000000000000110111010000000;
			12'b100010100100 		: log = 32'b00000000000000000110111010001010;
			12'b100010100101 		: log = 32'b00000000000000000110111010010101;
			12'b100010100110 		: log = 32'b00000000000000000110111010011111;
			12'b100010100111 		: log = 32'b00000000000000000110111010101010;
			12'b100010101000 		: log = 32'b00000000000000000110111010110100;
			12'b100010101001 		: log = 32'b00000000000000000110111010111110;
			12'b100010101010 		: log = 32'b00000000000000000110111011001001;
			12'b100010101011 		: log = 32'b00000000000000000110111011010011;
			12'b100010101100 		: log = 32'b00000000000000000110111011011110;
			12'b100010101101 		: log = 32'b00000000000000000110111011101000;
			12'b100010101110 		: log = 32'b00000000000000000110111011110010;
			12'b100010101111 		: log = 32'b00000000000000000110111011111101;
			12'b100010110000 		: log = 32'b00000000000000000110111100000111;
			12'b100010110001 		: log = 32'b00000000000000000110111100010001;
			12'b100010110010 		: log = 32'b00000000000000000110111100011100;
			12'b100010110011 		: log = 32'b00000000000000000110111100100110;
			12'b100010110100 		: log = 32'b00000000000000000110111100110000;
			12'b100010110101 		: log = 32'b00000000000000000110111100111011;
			12'b100010110110 		: log = 32'b00000000000000000110111101000101;
			12'b100010110111 		: log = 32'b00000000000000000110111101010000;
			12'b100010111000 		: log = 32'b00000000000000000110111101011010;
			12'b100010111001 		: log = 32'b00000000000000000110111101100100;
			12'b100010111010 		: log = 32'b00000000000000000110111101101111;
			12'b100010111011 		: log = 32'b00000000000000000110111101111001;
			12'b100010111100 		: log = 32'b00000000000000000110111110000011;
			12'b100010111101 		: log = 32'b00000000000000000110111110001110;
			12'b100010111110 		: log = 32'b00000000000000000110111110011000;
			12'b100010111111 		: log = 32'b00000000000000000110111110100010;
			12'b100011000000 		: log = 32'b00000000000000000110111110101101;
			12'b100011000001 		: log = 32'b00000000000000000110111110110111;
			12'b100011000010 		: log = 32'b00000000000000000110111111000001;
			12'b100011000011 		: log = 32'b00000000000000000110111111001100;
			12'b100011000100 		: log = 32'b00000000000000000110111111010110;
			12'b100011000101 		: log = 32'b00000000000000000110111111100000;
			12'b100011000110 		: log = 32'b00000000000000000110111111101011;
			12'b100011000111 		: log = 32'b00000000000000000110111111110101;
			12'b100011001000 		: log = 32'b00000000000000000110111111111111;
			12'b100011001001 		: log = 32'b00000000000000000111000000001010;
			12'b100011001010 		: log = 32'b00000000000000000111000000010100;
			12'b100011001011 		: log = 32'b00000000000000000111000000011110;
			12'b100011001100 		: log = 32'b00000000000000000111000000101001;
			12'b100011001101 		: log = 32'b00000000000000000111000000110011;
			12'b100011001110 		: log = 32'b00000000000000000111000000111101;
			12'b100011001111 		: log = 32'b00000000000000000111000001001000;
			12'b100011010000 		: log = 32'b00000000000000000111000001010010;
			12'b100011010001 		: log = 32'b00000000000000000111000001011100;
			12'b100011010010 		: log = 32'b00000000000000000111000001100111;
			12'b100011010011 		: log = 32'b00000000000000000111000001110001;
			12'b100011010100 		: log = 32'b00000000000000000111000001111011;
			12'b100011010101 		: log = 32'b00000000000000000111000010000110;
			12'b100011010110 		: log = 32'b00000000000000000111000010010000;
			12'b100011010111 		: log = 32'b00000000000000000111000010011010;
			12'b100011011000 		: log = 32'b00000000000000000111000010100100;
			12'b100011011001 		: log = 32'b00000000000000000111000010101111;
			12'b100011011010 		: log = 32'b00000000000000000111000010111001;
			12'b100011011011 		: log = 32'b00000000000000000111000011000011;
			12'b100011011100 		: log = 32'b00000000000000000111000011001110;
			12'b100011011101 		: log = 32'b00000000000000000111000011011000;
			12'b100011011110 		: log = 32'b00000000000000000111000011100010;
			12'b100011011111 		: log = 32'b00000000000000000111000011101101;
			12'b100011100000 		: log = 32'b00000000000000000111000011110111;
			12'b100011100001 		: log = 32'b00000000000000000111000100000001;
			12'b100011100010 		: log = 32'b00000000000000000111000100001011;
			12'b100011100011 		: log = 32'b00000000000000000111000100010110;
			12'b100011100100 		: log = 32'b00000000000000000111000100100000;
			12'b100011100101 		: log = 32'b00000000000000000111000100101010;
			12'b100011100110 		: log = 32'b00000000000000000111000100110101;
			12'b100011100111 		: log = 32'b00000000000000000111000100111111;
			12'b100011101000 		: log = 32'b00000000000000000111000101001001;
			12'b100011101001 		: log = 32'b00000000000000000111000101010011;
			12'b100011101010 		: log = 32'b00000000000000000111000101011110;
			12'b100011101011 		: log = 32'b00000000000000000111000101101000;
			12'b100011101100 		: log = 32'b00000000000000000111000101110010;
			12'b100011101101 		: log = 32'b00000000000000000111000101111101;
			12'b100011101110 		: log = 32'b00000000000000000111000110000111;
			12'b100011101111 		: log = 32'b00000000000000000111000110010001;
			12'b100011110000 		: log = 32'b00000000000000000111000110011011;
			12'b100011110001 		: log = 32'b00000000000000000111000110100110;
			12'b100011110010 		: log = 32'b00000000000000000111000110110000;
			12'b100011110011 		: log = 32'b00000000000000000111000110111010;
			12'b100011110100 		: log = 32'b00000000000000000111000111000100;
			12'b100011110101 		: log = 32'b00000000000000000111000111001111;
			12'b100011110110 		: log = 32'b00000000000000000111000111011001;
			12'b100011110111 		: log = 32'b00000000000000000111000111100011;
			12'b100011111000 		: log = 32'b00000000000000000111000111101101;
			12'b100011111001 		: log = 32'b00000000000000000111000111111000;
			12'b100011111010 		: log = 32'b00000000000000000111001000000010;
			12'b100011111011 		: log = 32'b00000000000000000111001000001100;
			12'b100011111100 		: log = 32'b00000000000000000111001000010110;
			12'b100011111101 		: log = 32'b00000000000000000111001000100001;
			12'b100011111110 		: log = 32'b00000000000000000111001000101011;
			12'b100011111111 		: log = 32'b00000000000000000111001000110101;
			12'b100100000000 		: log = 32'b00000000000000000111001000111111;
			12'b100100000001 		: log = 32'b00000000000000000111001001001010;
			12'b100100000010 		: log = 32'b00000000000000000111001001010100;
			12'b100100000011 		: log = 32'b00000000000000000111001001011110;
			12'b100100000100 		: log = 32'b00000000000000000111001001101000;
			12'b100100000101 		: log = 32'b00000000000000000111001001110011;
			12'b100100000110 		: log = 32'b00000000000000000111001001111101;
			12'b100100000111 		: log = 32'b00000000000000000111001010000111;
			12'b100100001000 		: log = 32'b00000000000000000111001010010001;
			12'b100100001001 		: log = 32'b00000000000000000111001010011011;
			12'b100100001010 		: log = 32'b00000000000000000111001010100110;
			12'b100100001011 		: log = 32'b00000000000000000111001010110000;
			12'b100100001100 		: log = 32'b00000000000000000111001010111010;
			12'b100100001101 		: log = 32'b00000000000000000111001011000100;
			12'b100100001110 		: log = 32'b00000000000000000111001011001111;
			12'b100100001111 		: log = 32'b00000000000000000111001011011001;
			12'b100100010000 		: log = 32'b00000000000000000111001011100011;
			12'b100100010001 		: log = 32'b00000000000000000111001011101101;
			12'b100100010010 		: log = 32'b00000000000000000111001011110111;
			12'b100100010011 		: log = 32'b00000000000000000111001100000010;
			12'b100100010100 		: log = 32'b00000000000000000111001100001100;
			12'b100100010101 		: log = 32'b00000000000000000111001100010110;
			12'b100100010110 		: log = 32'b00000000000000000111001100100000;
			12'b100100010111 		: log = 32'b00000000000000000111001100101010;
			12'b100100011000 		: log = 32'b00000000000000000111001100110101;
			12'b100100011001 		: log = 32'b00000000000000000111001100111111;
			12'b100100011010 		: log = 32'b00000000000000000111001101001001;
			12'b100100011011 		: log = 32'b00000000000000000111001101010011;
			12'b100100011100 		: log = 32'b00000000000000000111001101011101;
			12'b100100011101 		: log = 32'b00000000000000000111001101101000;
			12'b100100011110 		: log = 32'b00000000000000000111001101110010;
			12'b100100011111 		: log = 32'b00000000000000000111001101111100;
			12'b100100100000 		: log = 32'b00000000000000000111001110000110;
			12'b100100100001 		: log = 32'b00000000000000000111001110010000;
			12'b100100100010 		: log = 32'b00000000000000000111001110011011;
			12'b100100100011 		: log = 32'b00000000000000000111001110100101;
			12'b100100100100 		: log = 32'b00000000000000000111001110101111;
			12'b100100100101 		: log = 32'b00000000000000000111001110111001;
			12'b100100100110 		: log = 32'b00000000000000000111001111000011;
			12'b100100100111 		: log = 32'b00000000000000000111001111001110;
			12'b100100101000 		: log = 32'b00000000000000000111001111011000;
			12'b100100101001 		: log = 32'b00000000000000000111001111100010;
			12'b100100101010 		: log = 32'b00000000000000000111001111101100;
			12'b100100101011 		: log = 32'b00000000000000000111001111110110;
			12'b100100101100 		: log = 32'b00000000000000000111010000000000;
			12'b100100101101 		: log = 32'b00000000000000000111010000001011;
			12'b100100101110 		: log = 32'b00000000000000000111010000010101;
			12'b100100101111 		: log = 32'b00000000000000000111010000011111;
			12'b100100110000 		: log = 32'b00000000000000000111010000101001;
			12'b100100110001 		: log = 32'b00000000000000000111010000110011;
			12'b100100110010 		: log = 32'b00000000000000000111010000111101;
			12'b100100110011 		: log = 32'b00000000000000000111010001001000;
			12'b100100110100 		: log = 32'b00000000000000000111010001010010;
			12'b100100110101 		: log = 32'b00000000000000000111010001011100;
			12'b100100110110 		: log = 32'b00000000000000000111010001100110;
			12'b100100110111 		: log = 32'b00000000000000000111010001110000;
			12'b100100111000 		: log = 32'b00000000000000000111010001111010;
			12'b100100111001 		: log = 32'b00000000000000000111010010000100;
			12'b100100111010 		: log = 32'b00000000000000000111010010001111;
			12'b100100111011 		: log = 32'b00000000000000000111010010011001;
			12'b100100111100 		: log = 32'b00000000000000000111010010100011;
			12'b100100111101 		: log = 32'b00000000000000000111010010101101;
			12'b100100111110 		: log = 32'b00000000000000000111010010110111;
			12'b100100111111 		: log = 32'b00000000000000000111010011000001;
			12'b100101000000 		: log = 32'b00000000000000000111010011001011;
			12'b100101000001 		: log = 32'b00000000000000000111010011010110;
			12'b100101000010 		: log = 32'b00000000000000000111010011100000;
			12'b100101000011 		: log = 32'b00000000000000000111010011101010;
			12'b100101000100 		: log = 32'b00000000000000000111010011110100;
			12'b100101000101 		: log = 32'b00000000000000000111010011111110;
			12'b100101000110 		: log = 32'b00000000000000000111010100001000;
			12'b100101000111 		: log = 32'b00000000000000000111010100010010;
			12'b100101001000 		: log = 32'b00000000000000000111010100011101;
			12'b100101001001 		: log = 32'b00000000000000000111010100100111;
			12'b100101001010 		: log = 32'b00000000000000000111010100110001;
			12'b100101001011 		: log = 32'b00000000000000000111010100111011;
			12'b100101001100 		: log = 32'b00000000000000000111010101000101;
			12'b100101001101 		: log = 32'b00000000000000000111010101001111;
			12'b100101001110 		: log = 32'b00000000000000000111010101011001;
			12'b100101001111 		: log = 32'b00000000000000000111010101100011;
			12'b100101010000 		: log = 32'b00000000000000000111010101101101;
			12'b100101010001 		: log = 32'b00000000000000000111010101111000;
			12'b100101010010 		: log = 32'b00000000000000000111010110000010;
			12'b100101010011 		: log = 32'b00000000000000000111010110001100;
			12'b100101010100 		: log = 32'b00000000000000000111010110010110;
			12'b100101010101 		: log = 32'b00000000000000000111010110100000;
			12'b100101010110 		: log = 32'b00000000000000000111010110101010;
			12'b100101010111 		: log = 32'b00000000000000000111010110110100;
			12'b100101011000 		: log = 32'b00000000000000000111010110111110;
			12'b100101011001 		: log = 32'b00000000000000000111010111001000;
			12'b100101011010 		: log = 32'b00000000000000000111010111010011;
			12'b100101011011 		: log = 32'b00000000000000000111010111011101;
			12'b100101011100 		: log = 32'b00000000000000000111010111100111;
			12'b100101011101 		: log = 32'b00000000000000000111010111110001;
			12'b100101011110 		: log = 32'b00000000000000000111010111111011;
			12'b100101011111 		: log = 32'b00000000000000000111011000000101;
			12'b100101100000 		: log = 32'b00000000000000000111011000001111;
			12'b100101100001 		: log = 32'b00000000000000000111011000011001;
			12'b100101100010 		: log = 32'b00000000000000000111011000100011;
			12'b100101100011 		: log = 32'b00000000000000000111011000101101;
			12'b100101100100 		: log = 32'b00000000000000000111011000110111;
			12'b100101100101 		: log = 32'b00000000000000000111011001000010;
			12'b100101100110 		: log = 32'b00000000000000000111011001001100;
			12'b100101100111 		: log = 32'b00000000000000000111011001010110;
			12'b100101101000 		: log = 32'b00000000000000000111011001100000;
			12'b100101101001 		: log = 32'b00000000000000000111011001101010;
			12'b100101101010 		: log = 32'b00000000000000000111011001110100;
			12'b100101101011 		: log = 32'b00000000000000000111011001111110;
			12'b100101101100 		: log = 32'b00000000000000000111011010001000;
			12'b100101101101 		: log = 32'b00000000000000000111011010010010;
			12'b100101101110 		: log = 32'b00000000000000000111011010011100;
			12'b100101101111 		: log = 32'b00000000000000000111011010100110;
			12'b100101110000 		: log = 32'b00000000000000000111011010110000;
			12'b100101110001 		: log = 32'b00000000000000000111011010111010;
			12'b100101110010 		: log = 32'b00000000000000000111011011000100;
			12'b100101110011 		: log = 32'b00000000000000000111011011001111;
			12'b100101110100 		: log = 32'b00000000000000000111011011011001;
			12'b100101110101 		: log = 32'b00000000000000000111011011100011;
			12'b100101110110 		: log = 32'b00000000000000000111011011101101;
			12'b100101110111 		: log = 32'b00000000000000000111011011110111;
			12'b100101111000 		: log = 32'b00000000000000000111011100000001;
			12'b100101111001 		: log = 32'b00000000000000000111011100001011;
			12'b100101111010 		: log = 32'b00000000000000000111011100010101;
			12'b100101111011 		: log = 32'b00000000000000000111011100011111;
			12'b100101111100 		: log = 32'b00000000000000000111011100101001;
			12'b100101111101 		: log = 32'b00000000000000000111011100110011;
			12'b100101111110 		: log = 32'b00000000000000000111011100111101;
			12'b100101111111 		: log = 32'b00000000000000000111011101000111;
			12'b100110000000 		: log = 32'b00000000000000000111011101010001;
			12'b100110000001 		: log = 32'b00000000000000000111011101011011;
			12'b100110000010 		: log = 32'b00000000000000000111011101100101;
			12'b100110000011 		: log = 32'b00000000000000000111011101101111;
			12'b100110000100 		: log = 32'b00000000000000000111011101111001;
			12'b100110000101 		: log = 32'b00000000000000000111011110000011;
			12'b100110000110 		: log = 32'b00000000000000000111011110001101;
			12'b100110000111 		: log = 32'b00000000000000000111011110010111;
			12'b100110001000 		: log = 32'b00000000000000000111011110100001;
			12'b100110001001 		: log = 32'b00000000000000000111011110101011;
			12'b100110001010 		: log = 32'b00000000000000000111011110110101;
			12'b100110001011 		: log = 32'b00000000000000000111011110111111;
			12'b100110001100 		: log = 32'b00000000000000000111011111001010;
			12'b100110001101 		: log = 32'b00000000000000000111011111010100;
			12'b100110001110 		: log = 32'b00000000000000000111011111011110;
			12'b100110001111 		: log = 32'b00000000000000000111011111101000;
			12'b100110010000 		: log = 32'b00000000000000000111011111110010;
			12'b100110010001 		: log = 32'b00000000000000000111011111111100;
			12'b100110010010 		: log = 32'b00000000000000000111100000000110;
			12'b100110010011 		: log = 32'b00000000000000000111100000010000;
			12'b100110010100 		: log = 32'b00000000000000000111100000011010;
			12'b100110010101 		: log = 32'b00000000000000000111100000100100;
			12'b100110010110 		: log = 32'b00000000000000000111100000101110;
			12'b100110010111 		: log = 32'b00000000000000000111100000111000;
			12'b100110011000 		: log = 32'b00000000000000000111100001000010;
			12'b100110011001 		: log = 32'b00000000000000000111100001001100;
			12'b100110011010 		: log = 32'b00000000000000000111100001010110;
			12'b100110011011 		: log = 32'b00000000000000000111100001100000;
			12'b100110011100 		: log = 32'b00000000000000000111100001101010;
			12'b100110011101 		: log = 32'b00000000000000000111100001110100;
			12'b100110011110 		: log = 32'b00000000000000000111100001111110;
			12'b100110011111 		: log = 32'b00000000000000000111100010001000;
			12'b100110100000 		: log = 32'b00000000000000000111100010010010;
			12'b100110100001 		: log = 32'b00000000000000000111100010011100;
			12'b100110100010 		: log = 32'b00000000000000000111100010100110;
			12'b100110100011 		: log = 32'b00000000000000000111100010110000;
			12'b100110100100 		: log = 32'b00000000000000000111100010111010;
			12'b100110100101 		: log = 32'b00000000000000000111100011000100;
			12'b100110100110 		: log = 32'b00000000000000000111100011001110;
			12'b100110100111 		: log = 32'b00000000000000000111100011011000;
			12'b100110101000 		: log = 32'b00000000000000000111100011100001;
			12'b100110101001 		: log = 32'b00000000000000000111100011101011;
			12'b100110101010 		: log = 32'b00000000000000000111100011110101;
			12'b100110101011 		: log = 32'b00000000000000000111100011111111;
			12'b100110101100 		: log = 32'b00000000000000000111100100001001;
			12'b100110101101 		: log = 32'b00000000000000000111100100010011;
			12'b100110101110 		: log = 32'b00000000000000000111100100011101;
			12'b100110101111 		: log = 32'b00000000000000000111100100100111;
			12'b100110110000 		: log = 32'b00000000000000000111100100110001;
			12'b100110110001 		: log = 32'b00000000000000000111100100111011;
			12'b100110110010 		: log = 32'b00000000000000000111100101000101;
			12'b100110110011 		: log = 32'b00000000000000000111100101001111;
			12'b100110110100 		: log = 32'b00000000000000000111100101011001;
			12'b100110110101 		: log = 32'b00000000000000000111100101100011;
			12'b100110110110 		: log = 32'b00000000000000000111100101101101;
			12'b100110110111 		: log = 32'b00000000000000000111100101110111;
			12'b100110111000 		: log = 32'b00000000000000000111100110000001;
			12'b100110111001 		: log = 32'b00000000000000000111100110001011;
			12'b100110111010 		: log = 32'b00000000000000000111100110010101;
			12'b100110111011 		: log = 32'b00000000000000000111100110011111;
			12'b100110111100 		: log = 32'b00000000000000000111100110101001;
			12'b100110111101 		: log = 32'b00000000000000000111100110110011;
			12'b100110111110 		: log = 32'b00000000000000000111100110111101;
			12'b100110111111 		: log = 32'b00000000000000000111100111000111;
			12'b100111000000 		: log = 32'b00000000000000000111100111010001;
			12'b100111000001 		: log = 32'b00000000000000000111100111011010;
			12'b100111000010 		: log = 32'b00000000000000000111100111100100;
			12'b100111000011 		: log = 32'b00000000000000000111100111101110;
			12'b100111000100 		: log = 32'b00000000000000000111100111111000;
			12'b100111000101 		: log = 32'b00000000000000000111101000000010;
			12'b100111000110 		: log = 32'b00000000000000000111101000001100;
			12'b100111000111 		: log = 32'b00000000000000000111101000010110;
			12'b100111001000 		: log = 32'b00000000000000000111101000100000;
			12'b100111001001 		: log = 32'b00000000000000000111101000101010;
			12'b100111001010 		: log = 32'b00000000000000000111101000110100;
			12'b100111001011 		: log = 32'b00000000000000000111101000111110;
			12'b100111001100 		: log = 32'b00000000000000000111101001001000;
			12'b100111001101 		: log = 32'b00000000000000000111101001010010;
			12'b100111001110 		: log = 32'b00000000000000000111101001011100;
			12'b100111001111 		: log = 32'b00000000000000000111101001100101;
			12'b100111010000 		: log = 32'b00000000000000000111101001101111;
			12'b100111010001 		: log = 32'b00000000000000000111101001111001;
			12'b100111010010 		: log = 32'b00000000000000000111101010000011;
			12'b100111010011 		: log = 32'b00000000000000000111101010001101;
			12'b100111010100 		: log = 32'b00000000000000000111101010010111;
			12'b100111010101 		: log = 32'b00000000000000000111101010100001;
			12'b100111010110 		: log = 32'b00000000000000000111101010101011;
			12'b100111010111 		: log = 32'b00000000000000000111101010110101;
			12'b100111011000 		: log = 32'b00000000000000000111101010111111;
			12'b100111011001 		: log = 32'b00000000000000000111101011001001;
			12'b100111011010 		: log = 32'b00000000000000000111101011010011;
			12'b100111011011 		: log = 32'b00000000000000000111101011011100;
			12'b100111011100 		: log = 32'b00000000000000000111101011100110;
			12'b100111011101 		: log = 32'b00000000000000000111101011110000;
			12'b100111011110 		: log = 32'b00000000000000000111101011111010;
			12'b100111011111 		: log = 32'b00000000000000000111101100000100;
			12'b100111100000 		: log = 32'b00000000000000000111101100001110;
			12'b100111100001 		: log = 32'b00000000000000000111101100011000;
			12'b100111100010 		: log = 32'b00000000000000000111101100100010;
			12'b100111100011 		: log = 32'b00000000000000000111101100101100;
			12'b100111100100 		: log = 32'b00000000000000000111101100110101;
			12'b100111100101 		: log = 32'b00000000000000000111101100111111;
			12'b100111100110 		: log = 32'b00000000000000000111101101001001;
			12'b100111100111 		: log = 32'b00000000000000000111101101010011;
			12'b100111101000 		: log = 32'b00000000000000000111101101011101;
			12'b100111101001 		: log = 32'b00000000000000000111101101100111;
			12'b100111101010 		: log = 32'b00000000000000000111101101110001;
			12'b100111101011 		: log = 32'b00000000000000000111101101111011;
			12'b100111101100 		: log = 32'b00000000000000000111101110000101;
			12'b100111101101 		: log = 32'b00000000000000000111101110001110;
			12'b100111101110 		: log = 32'b00000000000000000111101110011000;
			12'b100111101111 		: log = 32'b00000000000000000111101110100010;
			12'b100111110000 		: log = 32'b00000000000000000111101110101100;
			12'b100111110001 		: log = 32'b00000000000000000111101110110110;
			12'b100111110010 		: log = 32'b00000000000000000111101111000000;
			12'b100111110011 		: log = 32'b00000000000000000111101111001010;
			12'b100111110100 		: log = 32'b00000000000000000111101111010011;
			12'b100111110101 		: log = 32'b00000000000000000111101111011101;
			12'b100111110110 		: log = 32'b00000000000000000111101111100111;
			12'b100111110111 		: log = 32'b00000000000000000111101111110001;
			12'b100111111000 		: log = 32'b00000000000000000111101111111011;
			12'b100111111001 		: log = 32'b00000000000000000111110000000101;
			12'b100111111010 		: log = 32'b00000000000000000111110000001111;
			12'b100111111011 		: log = 32'b00000000000000000111110000011000;
			12'b100111111100 		: log = 32'b00000000000000000111110000100010;
			12'b100111111101 		: log = 32'b00000000000000000111110000101100;
			12'b100111111110 		: log = 32'b00000000000000000111110000110110;
			12'b100111111111 		: log = 32'b00000000000000000111110001000000;
			12'b101000000000 		: log = 32'b00000000000000000111110001001010;
			12'b101000000001 		: log = 32'b00000000000000000111110001010100;
			12'b101000000010 		: log = 32'b00000000000000000111110001011101;
			12'b101000000011 		: log = 32'b00000000000000000111110001100111;
			12'b101000000100 		: log = 32'b00000000000000000111110001110001;
			12'b101000000101 		: log = 32'b00000000000000000111110001111011;
			12'b101000000110 		: log = 32'b00000000000000000111110010000101;
			12'b101000000111 		: log = 32'b00000000000000000111110010001111;
			12'b101000001000 		: log = 32'b00000000000000000111110010011000;
			12'b101000001001 		: log = 32'b00000000000000000111110010100010;
			12'b101000001010 		: log = 32'b00000000000000000111110010101100;
			12'b101000001011 		: log = 32'b00000000000000000111110010110110;
			12'b101000001100 		: log = 32'b00000000000000000111110011000000;
			12'b101000001101 		: log = 32'b00000000000000000111110011001010;
			12'b101000001110 		: log = 32'b00000000000000000111110011010011;
			12'b101000001111 		: log = 32'b00000000000000000111110011011101;
			12'b101000010000 		: log = 32'b00000000000000000111110011100111;
			12'b101000010001 		: log = 32'b00000000000000000111110011110001;
			12'b101000010010 		: log = 32'b00000000000000000111110011111011;
			12'b101000010011 		: log = 32'b00000000000000000111110100000101;
			12'b101000010100 		: log = 32'b00000000000000000111110100001110;
			12'b101000010101 		: log = 32'b00000000000000000111110100011000;
			12'b101000010110 		: log = 32'b00000000000000000111110100100010;
			12'b101000010111 		: log = 32'b00000000000000000111110100101100;
			12'b101000011000 		: log = 32'b00000000000000000111110100110110;
			12'b101000011001 		: log = 32'b00000000000000000111110100111111;
			12'b101000011010 		: log = 32'b00000000000000000111110101001001;
			12'b101000011011 		: log = 32'b00000000000000000111110101010011;
			12'b101000011100 		: log = 32'b00000000000000000111110101011101;
			12'b101000011101 		: log = 32'b00000000000000000111110101100111;
			12'b101000011110 		: log = 32'b00000000000000000111110101110000;
			12'b101000011111 		: log = 32'b00000000000000000111110101111010;
			12'b101000100000 		: log = 32'b00000000000000000111110110000100;
			12'b101000100001 		: log = 32'b00000000000000000111110110001110;
			12'b101000100010 		: log = 32'b00000000000000000111110110011000;
			12'b101000100011 		: log = 32'b00000000000000000111110110100001;
			12'b101000100100 		: log = 32'b00000000000000000111110110101011;
			12'b101000100101 		: log = 32'b00000000000000000111110110110101;
			12'b101000100110 		: log = 32'b00000000000000000111110110111111;
			12'b101000100111 		: log = 32'b00000000000000000111110111001001;
			12'b101000101000 		: log = 32'b00000000000000000111110111010010;
			12'b101000101001 		: log = 32'b00000000000000000111110111011100;
			12'b101000101010 		: log = 32'b00000000000000000111110111100110;
			12'b101000101011 		: log = 32'b00000000000000000111110111110000;
			12'b101000101100 		: log = 32'b00000000000000000111110111111010;
			12'b101000101101 		: log = 32'b00000000000000000111111000000011;
			12'b101000101110 		: log = 32'b00000000000000000111111000001101;
			12'b101000101111 		: log = 32'b00000000000000000111111000010111;
			12'b101000110000 		: log = 32'b00000000000000000111111000100001;
			12'b101000110001 		: log = 32'b00000000000000000111111000101010;
			12'b101000110010 		: log = 32'b00000000000000000111111000110100;
			12'b101000110011 		: log = 32'b00000000000000000111111000111110;
			12'b101000110100 		: log = 32'b00000000000000000111111001001000;
			12'b101000110101 		: log = 32'b00000000000000000111111001010010;
			12'b101000110110 		: log = 32'b00000000000000000111111001011011;
			12'b101000110111 		: log = 32'b00000000000000000111111001100101;
			12'b101000111000 		: log = 32'b00000000000000000111111001101111;
			12'b101000111001 		: log = 32'b00000000000000000111111001111001;
			12'b101000111010 		: log = 32'b00000000000000000111111010000010;
			12'b101000111011 		: log = 32'b00000000000000000111111010001100;
			12'b101000111100 		: log = 32'b00000000000000000111111010010110;
			12'b101000111101 		: log = 32'b00000000000000000111111010100000;
			12'b101000111110 		: log = 32'b00000000000000000111111010101001;
			12'b101000111111 		: log = 32'b00000000000000000111111010110011;
			12'b101001000000 		: log = 32'b00000000000000000111111010111101;
			12'b101001000001 		: log = 32'b00000000000000000111111011000111;
			12'b101001000010 		: log = 32'b00000000000000000111111011010000;
			12'b101001000011 		: log = 32'b00000000000000000111111011011010;
			12'b101001000100 		: log = 32'b00000000000000000111111011100100;
			12'b101001000101 		: log = 32'b00000000000000000111111011101110;
			12'b101001000110 		: log = 32'b00000000000000000111111011110111;
			12'b101001000111 		: log = 32'b00000000000000000111111100000001;
			12'b101001001000 		: log = 32'b00000000000000000111111100001011;
			12'b101001001001 		: log = 32'b00000000000000000111111100010101;
			12'b101001001010 		: log = 32'b00000000000000000111111100011110;
			12'b101001001011 		: log = 32'b00000000000000000111111100101000;
			12'b101001001100 		: log = 32'b00000000000000000111111100110010;
			12'b101001001101 		: log = 32'b00000000000000000111111100111100;
			12'b101001001110 		: log = 32'b00000000000000000111111101000101;
			12'b101001001111 		: log = 32'b00000000000000000111111101001111;
			12'b101001010000 		: log = 32'b00000000000000000111111101011001;
			12'b101001010001 		: log = 32'b00000000000000000111111101100010;
			12'b101001010010 		: log = 32'b00000000000000000111111101101100;
			12'b101001010011 		: log = 32'b00000000000000000111111101110110;
			12'b101001010100 		: log = 32'b00000000000000000111111110000000;
			12'b101001010101 		: log = 32'b00000000000000000111111110001001;
			12'b101001010110 		: log = 32'b00000000000000000111111110010011;
			12'b101001010111 		: log = 32'b00000000000000000111111110011101;
			12'b101001011000 		: log = 32'b00000000000000000111111110100111;
			12'b101001011001 		: log = 32'b00000000000000000111111110110000;
			12'b101001011010 		: log = 32'b00000000000000000111111110111010;
			12'b101001011011 		: log = 32'b00000000000000000111111111000100;
			12'b101001011100 		: log = 32'b00000000000000000111111111001101;
			12'b101001011101 		: log = 32'b00000000000000000111111111010111;
			12'b101001011110 		: log = 32'b00000000000000000111111111100001;
			12'b101001011111 		: log = 32'b00000000000000000111111111101011;
			12'b101001100000 		: log = 32'b00000000000000000111111111110100;
			12'b101001100001 		: log = 32'b00000000000000000111111111111110;
			12'b101001100010 		: log = 32'b00000000000000001000000000001000;
			12'b101001100011 		: log = 32'b00000000000000001000000000010001;
			12'b101001100100 		: log = 32'b00000000000000001000000000011011;
			12'b101001100101 		: log = 32'b00000000000000001000000000100101;
			12'b101001100110 		: log = 32'b00000000000000001000000000101110;
			12'b101001100111 		: log = 32'b00000000000000001000000000111000;
			12'b101001101000 		: log = 32'b00000000000000001000000001000010;
			12'b101001101001 		: log = 32'b00000000000000001000000001001100;
			12'b101001101010 		: log = 32'b00000000000000001000000001010101;
			12'b101001101011 		: log = 32'b00000000000000001000000001011111;
			12'b101001101100 		: log = 32'b00000000000000001000000001101001;
			12'b101001101101 		: log = 32'b00000000000000001000000001110010;
			12'b101001101110 		: log = 32'b00000000000000001000000001111100;
			12'b101001101111 		: log = 32'b00000000000000001000000010000110;
			12'b101001110000 		: log = 32'b00000000000000001000000010001111;
			12'b101001110001 		: log = 32'b00000000000000001000000010011001;
			12'b101001110010 		: log = 32'b00000000000000001000000010100011;
			12'b101001110011 		: log = 32'b00000000000000001000000010101100;
			12'b101001110100 		: log = 32'b00000000000000001000000010110110;
			12'b101001110101 		: log = 32'b00000000000000001000000011000000;
			12'b101001110110 		: log = 32'b00000000000000001000000011001001;
			12'b101001110111 		: log = 32'b00000000000000001000000011010011;
			12'b101001111000 		: log = 32'b00000000000000001000000011011101;
			12'b101001111001 		: log = 32'b00000000000000001000000011100110;
			12'b101001111010 		: log = 32'b00000000000000001000000011110000;
			12'b101001111011 		: log = 32'b00000000000000001000000011111010;
			12'b101001111100 		: log = 32'b00000000000000001000000100000011;
			12'b101001111101 		: log = 32'b00000000000000001000000100001101;
			12'b101001111110 		: log = 32'b00000000000000001000000100010111;
			12'b101001111111 		: log = 32'b00000000000000001000000100100000;
			12'b101010000000 		: log = 32'b00000000000000001000000100101010;
			12'b101010000001 		: log = 32'b00000000000000001000000100110100;
			12'b101010000010 		: log = 32'b00000000000000001000000100111101;
			12'b101010000011 		: log = 32'b00000000000000001000000101000111;
			12'b101010000100 		: log = 32'b00000000000000001000000101010001;
			12'b101010000101 		: log = 32'b00000000000000001000000101011010;
			12'b101010000110 		: log = 32'b00000000000000001000000101100100;
			12'b101010000111 		: log = 32'b00000000000000001000000101101110;
			12'b101010001000 		: log = 32'b00000000000000001000000101110111;
			12'b101010001001 		: log = 32'b00000000000000001000000110000001;
			12'b101010001010 		: log = 32'b00000000000000001000000110001011;
			12'b101010001011 		: log = 32'b00000000000000001000000110010100;
			12'b101010001100 		: log = 32'b00000000000000001000000110011110;
			12'b101010001101 		: log = 32'b00000000000000001000000110101000;
			12'b101010001110 		: log = 32'b00000000000000001000000110110001;
			12'b101010001111 		: log = 32'b00000000000000001000000110111011;
			12'b101010010000 		: log = 32'b00000000000000001000000111000100;
			12'b101010010001 		: log = 32'b00000000000000001000000111001110;
			12'b101010010010 		: log = 32'b00000000000000001000000111011000;
			12'b101010010011 		: log = 32'b00000000000000001000000111100001;
			12'b101010010100 		: log = 32'b00000000000000001000000111101011;
			12'b101010010101 		: log = 32'b00000000000000001000000111110101;
			12'b101010010110 		: log = 32'b00000000000000001000000111111110;
			12'b101010010111 		: log = 32'b00000000000000001000001000001000;
			12'b101010011000 		: log = 32'b00000000000000001000001000010010;
			12'b101010011001 		: log = 32'b00000000000000001000001000011011;
			12'b101010011010 		: log = 32'b00000000000000001000001000100101;
			12'b101010011011 		: log = 32'b00000000000000001000001000101110;
			12'b101010011100 		: log = 32'b00000000000000001000001000111000;
			12'b101010011101 		: log = 32'b00000000000000001000001001000010;
			12'b101010011110 		: log = 32'b00000000000000001000001001001011;
			12'b101010011111 		: log = 32'b00000000000000001000001001010101;
			12'b101010100000 		: log = 32'b00000000000000001000001001011110;
			12'b101010100001 		: log = 32'b00000000000000001000001001101000;
			12'b101010100010 		: log = 32'b00000000000000001000001001110010;
			12'b101010100011 		: log = 32'b00000000000000001000001001111011;
			12'b101010100100 		: log = 32'b00000000000000001000001010000101;
			12'b101010100101 		: log = 32'b00000000000000001000001010001111;
			12'b101010100110 		: log = 32'b00000000000000001000001010011000;
			12'b101010100111 		: log = 32'b00000000000000001000001010100010;
			12'b101010101000 		: log = 32'b00000000000000001000001010101011;
			12'b101010101001 		: log = 32'b00000000000000001000001010110101;
			12'b101010101010 		: log = 32'b00000000000000001000001010111111;
			12'b101010101011 		: log = 32'b00000000000000001000001011001000;
			12'b101010101100 		: log = 32'b00000000000000001000001011010010;
			12'b101010101101 		: log = 32'b00000000000000001000001011011011;
			12'b101010101110 		: log = 32'b00000000000000001000001011100101;
			12'b101010101111 		: log = 32'b00000000000000001000001011101111;
			12'b101010110000 		: log = 32'b00000000000000001000001011111000;
			12'b101010110001 		: log = 32'b00000000000000001000001100000010;
			12'b101010110010 		: log = 32'b00000000000000001000001100001011;
			12'b101010110011 		: log = 32'b00000000000000001000001100010101;
			12'b101010110100 		: log = 32'b00000000000000001000001100011111;
			12'b101010110101 		: log = 32'b00000000000000001000001100101000;
			12'b101010110110 		: log = 32'b00000000000000001000001100110010;
			12'b101010110111 		: log = 32'b00000000000000001000001100111011;
			12'b101010111000 		: log = 32'b00000000000000001000001101000101;
			12'b101010111001 		: log = 32'b00000000000000001000001101001110;
			12'b101010111010 		: log = 32'b00000000000000001000001101011000;
			12'b101010111011 		: log = 32'b00000000000000001000001101100010;
			12'b101010111100 		: log = 32'b00000000000000001000001101101011;
			12'b101010111101 		: log = 32'b00000000000000001000001101110101;
			12'b101010111110 		: log = 32'b00000000000000001000001101111110;
			12'b101010111111 		: log = 32'b00000000000000001000001110001000;
			12'b101011000000 		: log = 32'b00000000000000001000001110010001;
			12'b101011000001 		: log = 32'b00000000000000001000001110011011;
			12'b101011000010 		: log = 32'b00000000000000001000001110100101;
			12'b101011000011 		: log = 32'b00000000000000001000001110101110;
			12'b101011000100 		: log = 32'b00000000000000001000001110111000;
			12'b101011000101 		: log = 32'b00000000000000001000001111000001;
			12'b101011000110 		: log = 32'b00000000000000001000001111001011;
			12'b101011000111 		: log = 32'b00000000000000001000001111010100;
			12'b101011001000 		: log = 32'b00000000000000001000001111011110;
			12'b101011001001 		: log = 32'b00000000000000001000001111101000;
			12'b101011001010 		: log = 32'b00000000000000001000001111110001;
			12'b101011001011 		: log = 32'b00000000000000001000001111111011;
			12'b101011001100 		: log = 32'b00000000000000001000010000000100;
			12'b101011001101 		: log = 32'b00000000000000001000010000001110;
			12'b101011001110 		: log = 32'b00000000000000001000010000010111;
			12'b101011001111 		: log = 32'b00000000000000001000010000100001;
			12'b101011010000 		: log = 32'b00000000000000001000010000101010;
			12'b101011010001 		: log = 32'b00000000000000001000010000110100;
			12'b101011010010 		: log = 32'b00000000000000001000010000111101;
			12'b101011010011 		: log = 32'b00000000000000001000010001000111;
			12'b101011010100 		: log = 32'b00000000000000001000010001010001;
			12'b101011010101 		: log = 32'b00000000000000001000010001011010;
			12'b101011010110 		: log = 32'b00000000000000001000010001100100;
			12'b101011010111 		: log = 32'b00000000000000001000010001101101;
			12'b101011011000 		: log = 32'b00000000000000001000010001110111;
			12'b101011011001 		: log = 32'b00000000000000001000010010000000;
			12'b101011011010 		: log = 32'b00000000000000001000010010001010;
			12'b101011011011 		: log = 32'b00000000000000001000010010010011;
			12'b101011011100 		: log = 32'b00000000000000001000010010011101;
			12'b101011011101 		: log = 32'b00000000000000001000010010100110;
			12'b101011011110 		: log = 32'b00000000000000001000010010110000;
			12'b101011011111 		: log = 32'b00000000000000001000010010111001;
			12'b101011100000 		: log = 32'b00000000000000001000010011000011;
			12'b101011100001 		: log = 32'b00000000000000001000010011001101;
			12'b101011100010 		: log = 32'b00000000000000001000010011010110;
			12'b101011100011 		: log = 32'b00000000000000001000010011100000;
			12'b101011100100 		: log = 32'b00000000000000001000010011101001;
			12'b101011100101 		: log = 32'b00000000000000001000010011110011;
			12'b101011100110 		: log = 32'b00000000000000001000010011111100;
			12'b101011100111 		: log = 32'b00000000000000001000010100000110;
			12'b101011101000 		: log = 32'b00000000000000001000010100001111;
			12'b101011101001 		: log = 32'b00000000000000001000010100011001;
			12'b101011101010 		: log = 32'b00000000000000001000010100100010;
			12'b101011101011 		: log = 32'b00000000000000001000010100101100;
			12'b101011101100 		: log = 32'b00000000000000001000010100110101;
			12'b101011101101 		: log = 32'b00000000000000001000010100111111;
			12'b101011101110 		: log = 32'b00000000000000001000010101001000;
			12'b101011101111 		: log = 32'b00000000000000001000010101010010;
			12'b101011110000 		: log = 32'b00000000000000001000010101011011;
			12'b101011110001 		: log = 32'b00000000000000001000010101100101;
			12'b101011110010 		: log = 32'b00000000000000001000010101101110;
			12'b101011110011 		: log = 32'b00000000000000001000010101111000;
			12'b101011110100 		: log = 32'b00000000000000001000010110000001;
			12'b101011110101 		: log = 32'b00000000000000001000010110001011;
			12'b101011110110 		: log = 32'b00000000000000001000010110010100;
			12'b101011110111 		: log = 32'b00000000000000001000010110011110;
			12'b101011111000 		: log = 32'b00000000000000001000010110100111;
			12'b101011111001 		: log = 32'b00000000000000001000010110110001;
			12'b101011111010 		: log = 32'b00000000000000001000010110111010;
			12'b101011111011 		: log = 32'b00000000000000001000010111000100;
			12'b101011111100 		: log = 32'b00000000000000001000010111001101;
			12'b101011111101 		: log = 32'b00000000000000001000010111010111;
			12'b101011111110 		: log = 32'b00000000000000001000010111100000;
			12'b101011111111 		: log = 32'b00000000000000001000010111101010;
			12'b101100000000 		: log = 32'b00000000000000001000010111110011;
			12'b101100000001 		: log = 32'b00000000000000001000010111111101;
			12'b101100000010 		: log = 32'b00000000000000001000011000000110;
			12'b101100000011 		: log = 32'b00000000000000001000011000010000;
			12'b101100000100 		: log = 32'b00000000000000001000011000011001;
			12'b101100000101 		: log = 32'b00000000000000001000011000100010;
			12'b101100000110 		: log = 32'b00000000000000001000011000101100;
			12'b101100000111 		: log = 32'b00000000000000001000011000110101;
			12'b101100001000 		: log = 32'b00000000000000001000011000111111;
			12'b101100001001 		: log = 32'b00000000000000001000011001001000;
			12'b101100001010 		: log = 32'b00000000000000001000011001010010;
			12'b101100001011 		: log = 32'b00000000000000001000011001011011;
			12'b101100001100 		: log = 32'b00000000000000001000011001100101;
			12'b101100001101 		: log = 32'b00000000000000001000011001101110;
			12'b101100001110 		: log = 32'b00000000000000001000011001111000;
			12'b101100001111 		: log = 32'b00000000000000001000011010000001;
			12'b101100010000 		: log = 32'b00000000000000001000011010001011;
			12'b101100010001 		: log = 32'b00000000000000001000011010010100;
			12'b101100010010 		: log = 32'b00000000000000001000011010011110;
			12'b101100010011 		: log = 32'b00000000000000001000011010100111;
			12'b101100010100 		: log = 32'b00000000000000001000011010110000;
			12'b101100010101 		: log = 32'b00000000000000001000011010111010;
			12'b101100010110 		: log = 32'b00000000000000001000011011000011;
			12'b101100010111 		: log = 32'b00000000000000001000011011001101;
			12'b101100011000 		: log = 32'b00000000000000001000011011010110;
			12'b101100011001 		: log = 32'b00000000000000001000011011100000;
			12'b101100011010 		: log = 32'b00000000000000001000011011101001;
			12'b101100011011 		: log = 32'b00000000000000001000011011110011;
			12'b101100011100 		: log = 32'b00000000000000001000011011111100;
			12'b101100011101 		: log = 32'b00000000000000001000011100000101;
			12'b101100011110 		: log = 32'b00000000000000001000011100001111;
			12'b101100011111 		: log = 32'b00000000000000001000011100011000;
			12'b101100100000 		: log = 32'b00000000000000001000011100100010;
			12'b101100100001 		: log = 32'b00000000000000001000011100101011;
			12'b101100100010 		: log = 32'b00000000000000001000011100110101;
			12'b101100100011 		: log = 32'b00000000000000001000011100111110;
			12'b101100100100 		: log = 32'b00000000000000001000011101001000;
			12'b101100100101 		: log = 32'b00000000000000001000011101010001;
			12'b101100100110 		: log = 32'b00000000000000001000011101011010;
			12'b101100100111 		: log = 32'b00000000000000001000011101100100;
			12'b101100101000 		: log = 32'b00000000000000001000011101101101;
			12'b101100101001 		: log = 32'b00000000000000001000011101110111;
			12'b101100101010 		: log = 32'b00000000000000001000011110000000;
			12'b101100101011 		: log = 32'b00000000000000001000011110001010;
			12'b101100101100 		: log = 32'b00000000000000001000011110010011;
			12'b101100101101 		: log = 32'b00000000000000001000011110011100;
			12'b101100101110 		: log = 32'b00000000000000001000011110100110;
			12'b101100101111 		: log = 32'b00000000000000001000011110101111;
			12'b101100110000 		: log = 32'b00000000000000001000011110111001;
			12'b101100110001 		: log = 32'b00000000000000001000011111000010;
			12'b101100110010 		: log = 32'b00000000000000001000011111001011;
			12'b101100110011 		: log = 32'b00000000000000001000011111010101;
			12'b101100110100 		: log = 32'b00000000000000001000011111011110;
			12'b101100110101 		: log = 32'b00000000000000001000011111101000;
			12'b101100110110 		: log = 32'b00000000000000001000011111110001;
			12'b101100110111 		: log = 32'b00000000000000001000011111111011;
			12'b101100111000 		: log = 32'b00000000000000001000100000000100;
			12'b101100111001 		: log = 32'b00000000000000001000100000001101;
			12'b101100111010 		: log = 32'b00000000000000001000100000010111;
			12'b101100111011 		: log = 32'b00000000000000001000100000100000;
			12'b101100111100 		: log = 32'b00000000000000001000100000101010;
			12'b101100111101 		: log = 32'b00000000000000001000100000110011;
			12'b101100111110 		: log = 32'b00000000000000001000100000111100;
			12'b101100111111 		: log = 32'b00000000000000001000100001000110;
			12'b101101000000 		: log = 32'b00000000000000001000100001001111;
			12'b101101000001 		: log = 32'b00000000000000001000100001011001;
			12'b101101000010 		: log = 32'b00000000000000001000100001100010;
			12'b101101000011 		: log = 32'b00000000000000001000100001101011;
			12'b101101000100 		: log = 32'b00000000000000001000100001110101;
			12'b101101000101 		: log = 32'b00000000000000001000100001111110;
			12'b101101000110 		: log = 32'b00000000000000001000100010000111;
			12'b101101000111 		: log = 32'b00000000000000001000100010010001;
			12'b101101001000 		: log = 32'b00000000000000001000100010011010;
			12'b101101001001 		: log = 32'b00000000000000001000100010100100;
			12'b101101001010 		: log = 32'b00000000000000001000100010101101;
			12'b101101001011 		: log = 32'b00000000000000001000100010110110;
			12'b101101001100 		: log = 32'b00000000000000001000100011000000;
			12'b101101001101 		: log = 32'b00000000000000001000100011001001;
			12'b101101001110 		: log = 32'b00000000000000001000100011010011;
			12'b101101001111 		: log = 32'b00000000000000001000100011011100;
			12'b101101010000 		: log = 32'b00000000000000001000100011100101;
			12'b101101010001 		: log = 32'b00000000000000001000100011101111;
			12'b101101010010 		: log = 32'b00000000000000001000100011111000;
			12'b101101010011 		: log = 32'b00000000000000001000100100000001;
			12'b101101010100 		: log = 32'b00000000000000001000100100001011;
			12'b101101010101 		: log = 32'b00000000000000001000100100010100;
			12'b101101010110 		: log = 32'b00000000000000001000100100011101;
			12'b101101010111 		: log = 32'b00000000000000001000100100100111;
			12'b101101011000 		: log = 32'b00000000000000001000100100110000;
			12'b101101011001 		: log = 32'b00000000000000001000100100111010;
			12'b101101011010 		: log = 32'b00000000000000001000100101000011;
			12'b101101011011 		: log = 32'b00000000000000001000100101001100;
			12'b101101011100 		: log = 32'b00000000000000001000100101010110;
			12'b101101011101 		: log = 32'b00000000000000001000100101011111;
			12'b101101011110 		: log = 32'b00000000000000001000100101101000;
			12'b101101011111 		: log = 32'b00000000000000001000100101110010;
			12'b101101100000 		: log = 32'b00000000000000001000100101111011;
			12'b101101100001 		: log = 32'b00000000000000001000100110000100;
			12'b101101100010 		: log = 32'b00000000000000001000100110001110;
			12'b101101100011 		: log = 32'b00000000000000001000100110010111;
			12'b101101100100 		: log = 32'b00000000000000001000100110100000;
			12'b101101100101 		: log = 32'b00000000000000001000100110101010;
			12'b101101100110 		: log = 32'b00000000000000001000100110110011;
			12'b101101100111 		: log = 32'b00000000000000001000100110111100;
			12'b101101101000 		: log = 32'b00000000000000001000100111000110;
			12'b101101101001 		: log = 32'b00000000000000001000100111001111;
			12'b101101101010 		: log = 32'b00000000000000001000100111011000;
			12'b101101101011 		: log = 32'b00000000000000001000100111100010;
			12'b101101101100 		: log = 32'b00000000000000001000100111101011;
			12'b101101101101 		: log = 32'b00000000000000001000100111110101;
			12'b101101101110 		: log = 32'b00000000000000001000100111111110;
			12'b101101101111 		: log = 32'b00000000000000001000101000000111;
			12'b101101110000 		: log = 32'b00000000000000001000101000010001;
			12'b101101110001 		: log = 32'b00000000000000001000101000011010;
			12'b101101110010 		: log = 32'b00000000000000001000101000100011;
			12'b101101110011 		: log = 32'b00000000000000001000101000101100;
			12'b101101110100 		: log = 32'b00000000000000001000101000110110;
			12'b101101110101 		: log = 32'b00000000000000001000101000111111;
			12'b101101110110 		: log = 32'b00000000000000001000101001001000;
			12'b101101110111 		: log = 32'b00000000000000001000101001010010;
			12'b101101111000 		: log = 32'b00000000000000001000101001011011;
			12'b101101111001 		: log = 32'b00000000000000001000101001100100;
			12'b101101111010 		: log = 32'b00000000000000001000101001101110;
			12'b101101111011 		: log = 32'b00000000000000001000101001110111;
			12'b101101111100 		: log = 32'b00000000000000001000101010000000;
			12'b101101111101 		: log = 32'b00000000000000001000101010001010;
			12'b101101111110 		: log = 32'b00000000000000001000101010010011;
			12'b101101111111 		: log = 32'b00000000000000001000101010011100;
			12'b101110000000 		: log = 32'b00000000000000001000101010100110;
			12'b101110000001 		: log = 32'b00000000000000001000101010101111;
			12'b101110000010 		: log = 32'b00000000000000001000101010111000;
			12'b101110000011 		: log = 32'b00000000000000001000101011000010;
			12'b101110000100 		: log = 32'b00000000000000001000101011001011;
			12'b101110000101 		: log = 32'b00000000000000001000101011010100;
			12'b101110000110 		: log = 32'b00000000000000001000101011011101;
			12'b101110000111 		: log = 32'b00000000000000001000101011100111;
			12'b101110001000 		: log = 32'b00000000000000001000101011110000;
			12'b101110001001 		: log = 32'b00000000000000001000101011111001;
			12'b101110001010 		: log = 32'b00000000000000001000101100000011;
			12'b101110001011 		: log = 32'b00000000000000001000101100001100;
			12'b101110001100 		: log = 32'b00000000000000001000101100010101;
			12'b101110001101 		: log = 32'b00000000000000001000101100011111;
			12'b101110001110 		: log = 32'b00000000000000001000101100101000;
			12'b101110001111 		: log = 32'b00000000000000001000101100110001;
			12'b101110010000 		: log = 32'b00000000000000001000101100111010;
			12'b101110010001 		: log = 32'b00000000000000001000101101000100;
			12'b101110010010 		: log = 32'b00000000000000001000101101001101;
			12'b101110010011 		: log = 32'b00000000000000001000101101010110;
			12'b101110010100 		: log = 32'b00000000000000001000101101100000;
			12'b101110010101 		: log = 32'b00000000000000001000101101101001;
			12'b101110010110 		: log = 32'b00000000000000001000101101110010;
			12'b101110010111 		: log = 32'b00000000000000001000101101111011;
			12'b101110011000 		: log = 32'b00000000000000001000101110000101;
			12'b101110011001 		: log = 32'b00000000000000001000101110001110;
			12'b101110011010 		: log = 32'b00000000000000001000101110010111;
			12'b101110011011 		: log = 32'b00000000000000001000101110100000;
			12'b101110011100 		: log = 32'b00000000000000001000101110101010;
			12'b101110011101 		: log = 32'b00000000000000001000101110110011;
			12'b101110011110 		: log = 32'b00000000000000001000101110111100;
			12'b101110011111 		: log = 32'b00000000000000001000101111000110;
			12'b101110100000 		: log = 32'b00000000000000001000101111001111;
			12'b101110100001 		: log = 32'b00000000000000001000101111011000;
			12'b101110100010 		: log = 32'b00000000000000001000101111100001;
			12'b101110100011 		: log = 32'b00000000000000001000101111101011;
			12'b101110100100 		: log = 32'b00000000000000001000101111110100;
			12'b101110100101 		: log = 32'b00000000000000001000101111111101;
			12'b101110100110 		: log = 32'b00000000000000001000110000000110;
			12'b101110100111 		: log = 32'b00000000000000001000110000010000;
			12'b101110101000 		: log = 32'b00000000000000001000110000011001;
			12'b101110101001 		: log = 32'b00000000000000001000110000100010;
			12'b101110101010 		: log = 32'b00000000000000001000110000101011;
			12'b101110101011 		: log = 32'b00000000000000001000110000110101;
			12'b101110101100 		: log = 32'b00000000000000001000110000111110;
			12'b101110101101 		: log = 32'b00000000000000001000110001000111;
			12'b101110101110 		: log = 32'b00000000000000001000110001010000;
			12'b101110101111 		: log = 32'b00000000000000001000110001011010;
			12'b101110110000 		: log = 32'b00000000000000001000110001100011;
			12'b101110110001 		: log = 32'b00000000000000001000110001101100;
			12'b101110110010 		: log = 32'b00000000000000001000110001110101;
			12'b101110110011 		: log = 32'b00000000000000001000110001111111;
			12'b101110110100 		: log = 32'b00000000000000001000110010001000;
			12'b101110110101 		: log = 32'b00000000000000001000110010010001;
			12'b101110110110 		: log = 32'b00000000000000001000110010011010;
			12'b101110110111 		: log = 32'b00000000000000001000110010100100;
			12'b101110111000 		: log = 32'b00000000000000001000110010101101;
			12'b101110111001 		: log = 32'b00000000000000001000110010110110;
			12'b101110111010 		: log = 32'b00000000000000001000110010111111;
			12'b101110111011 		: log = 32'b00000000000000001000110011001001;
			12'b101110111100 		: log = 32'b00000000000000001000110011010010;
			12'b101110111101 		: log = 32'b00000000000000001000110011011011;
			12'b101110111110 		: log = 32'b00000000000000001000110011100100;
			12'b101110111111 		: log = 32'b00000000000000001000110011101101;
			12'b101111000000 		: log = 32'b00000000000000001000110011110111;
			12'b101111000001 		: log = 32'b00000000000000001000110100000000;
			12'b101111000010 		: log = 32'b00000000000000001000110100001001;
			12'b101111000011 		: log = 32'b00000000000000001000110100010010;
			12'b101111000100 		: log = 32'b00000000000000001000110100011100;
			12'b101111000101 		: log = 32'b00000000000000001000110100100101;
			12'b101111000110 		: log = 32'b00000000000000001000110100101110;
			12'b101111000111 		: log = 32'b00000000000000001000110100110111;
			12'b101111001000 		: log = 32'b00000000000000001000110101000000;
			12'b101111001001 		: log = 32'b00000000000000001000110101001010;
			12'b101111001010 		: log = 32'b00000000000000001000110101010011;
			12'b101111001011 		: log = 32'b00000000000000001000110101011100;
			12'b101111001100 		: log = 32'b00000000000000001000110101100101;
			12'b101111001101 		: log = 32'b00000000000000001000110101101111;
			12'b101111001110 		: log = 32'b00000000000000001000110101111000;
			12'b101111001111 		: log = 32'b00000000000000001000110110000001;
			12'b101111010000 		: log = 32'b00000000000000001000110110001010;
			12'b101111010001 		: log = 32'b00000000000000001000110110010011;
			12'b101111010010 		: log = 32'b00000000000000001000110110011101;
			12'b101111010011 		: log = 32'b00000000000000001000110110100110;
			12'b101111010100 		: log = 32'b00000000000000001000110110101111;
			12'b101111010101 		: log = 32'b00000000000000001000110110111000;
			12'b101111010110 		: log = 32'b00000000000000001000110111000001;
			12'b101111010111 		: log = 32'b00000000000000001000110111001011;
			12'b101111011000 		: log = 32'b00000000000000001000110111010100;
			12'b101111011001 		: log = 32'b00000000000000001000110111011101;
			12'b101111011010 		: log = 32'b00000000000000001000110111100110;
			12'b101111011011 		: log = 32'b00000000000000001000110111101111;
			12'b101111011100 		: log = 32'b00000000000000001000110111111001;
			12'b101111011101 		: log = 32'b00000000000000001000111000000010;
			12'b101111011110 		: log = 32'b00000000000000001000111000001011;
			12'b101111011111 		: log = 32'b00000000000000001000111000010100;
			12'b101111100000 		: log = 32'b00000000000000001000111000011101;
			12'b101111100001 		: log = 32'b00000000000000001000111000100110;
			12'b101111100010 		: log = 32'b00000000000000001000111000110000;
			12'b101111100011 		: log = 32'b00000000000000001000111000111001;
			12'b101111100100 		: log = 32'b00000000000000001000111001000010;
			12'b101111100101 		: log = 32'b00000000000000001000111001001011;
			12'b101111100110 		: log = 32'b00000000000000001000111001010100;
			12'b101111100111 		: log = 32'b00000000000000001000111001011110;
			12'b101111101000 		: log = 32'b00000000000000001000111001100111;
			12'b101111101001 		: log = 32'b00000000000000001000111001110000;
			12'b101111101010 		: log = 32'b00000000000000001000111001111001;
			12'b101111101011 		: log = 32'b00000000000000001000111010000010;
			12'b101111101100 		: log = 32'b00000000000000001000111010001011;
			12'b101111101101 		: log = 32'b00000000000000001000111010010101;
			12'b101111101110 		: log = 32'b00000000000000001000111010011110;
			12'b101111101111 		: log = 32'b00000000000000001000111010100111;
			12'b101111110000 		: log = 32'b00000000000000001000111010110000;
			12'b101111110001 		: log = 32'b00000000000000001000111010111001;
			12'b101111110010 		: log = 32'b00000000000000001000111011000010;
			12'b101111110011 		: log = 32'b00000000000000001000111011001100;
			12'b101111110100 		: log = 32'b00000000000000001000111011010101;
			12'b101111110101 		: log = 32'b00000000000000001000111011011110;
			12'b101111110110 		: log = 32'b00000000000000001000111011100111;
			12'b101111110111 		: log = 32'b00000000000000001000111011110000;
			12'b101111111000 		: log = 32'b00000000000000001000111011111001;
			12'b101111111001 		: log = 32'b00000000000000001000111100000010;
			12'b101111111010 		: log = 32'b00000000000000001000111100001100;
			12'b101111111011 		: log = 32'b00000000000000001000111100010101;
			12'b101111111100 		: log = 32'b00000000000000001000111100011110;
			12'b101111111101 		: log = 32'b00000000000000001000111100100111;
			12'b101111111110 		: log = 32'b00000000000000001000111100110000;
			12'b101111111111 		: log = 32'b00000000000000001000111100111001;
			12'b110000000000 		: log = 32'b00000000000000001000111101000010;
			12'b110000000001 		: log = 32'b00000000000000001000111101001100;
			12'b110000000010 		: log = 32'b00000000000000001000111101010101;
			12'b110000000011 		: log = 32'b00000000000000001000111101011110;
			12'b110000000100 		: log = 32'b00000000000000001000111101100111;
			12'b110000000101 		: log = 32'b00000000000000001000111101110000;
			12'b110000000110 		: log = 32'b00000000000000001000111101111001;
			12'b110000000111 		: log = 32'b00000000000000001000111110000010;
			12'b110000001000 		: log = 32'b00000000000000001000111110001100;
			12'b110000001001 		: log = 32'b00000000000000001000111110010101;
			12'b110000001010 		: log = 32'b00000000000000001000111110011110;
			12'b110000001011 		: log = 32'b00000000000000001000111110100111;
			12'b110000001100 		: log = 32'b00000000000000001000111110110000;
			12'b110000001101 		: log = 32'b00000000000000001000111110111001;
			12'b110000001110 		: log = 32'b00000000000000001000111111000010;
			12'b110000001111 		: log = 32'b00000000000000001000111111001011;
			12'b110000010000 		: log = 32'b00000000000000001000111111010101;
			12'b110000010001 		: log = 32'b00000000000000001000111111011110;
			12'b110000010010 		: log = 32'b00000000000000001000111111100111;
			12'b110000010011 		: log = 32'b00000000000000001000111111110000;
			12'b110000010100 		: log = 32'b00000000000000001000111111111001;
			12'b110000010101 		: log = 32'b00000000000000001001000000000010;
			12'b110000010110 		: log = 32'b00000000000000001001000000001011;
			12'b110000010111 		: log = 32'b00000000000000001001000000010100;
			12'b110000011000 		: log = 32'b00000000000000001001000000011110;
			12'b110000011001 		: log = 32'b00000000000000001001000000100111;
			12'b110000011010 		: log = 32'b00000000000000001001000000110000;
			12'b110000011011 		: log = 32'b00000000000000001001000000111001;
			12'b110000011100 		: log = 32'b00000000000000001001000001000010;
			12'b110000011101 		: log = 32'b00000000000000001001000001001011;
			12'b110000011110 		: log = 32'b00000000000000001001000001010100;
			12'b110000011111 		: log = 32'b00000000000000001001000001011101;
			12'b110000100000 		: log = 32'b00000000000000001001000001100110;
			12'b110000100001 		: log = 32'b00000000000000001001000001110000;
			12'b110000100010 		: log = 32'b00000000000000001001000001111001;
			12'b110000100011 		: log = 32'b00000000000000001001000010000010;
			12'b110000100100 		: log = 32'b00000000000000001001000010001011;
			12'b110000100101 		: log = 32'b00000000000000001001000010010100;
			12'b110000100110 		: log = 32'b00000000000000001001000010011101;
			12'b110000100111 		: log = 32'b00000000000000001001000010100110;
			12'b110000101000 		: log = 32'b00000000000000001001000010101111;
			12'b110000101001 		: log = 32'b00000000000000001001000010111000;
			12'b110000101010 		: log = 32'b00000000000000001001000011000001;
			12'b110000101011 		: log = 32'b00000000000000001001000011001010;
			12'b110000101100 		: log = 32'b00000000000000001001000011010100;
			12'b110000101101 		: log = 32'b00000000000000001001000011011101;
			12'b110000101110 		: log = 32'b00000000000000001001000011100110;
			12'b110000101111 		: log = 32'b00000000000000001001000011101111;
			12'b110000110000 		: log = 32'b00000000000000001001000011111000;
			12'b110000110001 		: log = 32'b00000000000000001001000100000001;
			12'b110000110010 		: log = 32'b00000000000000001001000100001010;
			12'b110000110011 		: log = 32'b00000000000000001001000100010011;
			12'b110000110100 		: log = 32'b00000000000000001001000100011100;
			12'b110000110101 		: log = 32'b00000000000000001001000100100101;
			12'b110000110110 		: log = 32'b00000000000000001001000100101110;
			12'b110000110111 		: log = 32'b00000000000000001001000100110111;
			12'b110000111000 		: log = 32'b00000000000000001001000101000000;
			12'b110000111001 		: log = 32'b00000000000000001001000101001010;
			12'b110000111010 		: log = 32'b00000000000000001001000101010011;
			12'b110000111011 		: log = 32'b00000000000000001001000101011100;
			12'b110000111100 		: log = 32'b00000000000000001001000101100101;
			12'b110000111101 		: log = 32'b00000000000000001001000101101110;
			12'b110000111110 		: log = 32'b00000000000000001001000101110111;
			12'b110000111111 		: log = 32'b00000000000000001001000110000000;
			12'b110001000000 		: log = 32'b00000000000000001001000110001001;
			12'b110001000001 		: log = 32'b00000000000000001001000110010010;
			12'b110001000010 		: log = 32'b00000000000000001001000110011011;
			12'b110001000011 		: log = 32'b00000000000000001001000110100100;
			12'b110001000100 		: log = 32'b00000000000000001001000110101101;
			12'b110001000101 		: log = 32'b00000000000000001001000110110110;
			12'b110001000110 		: log = 32'b00000000000000001001000110111111;
			12'b110001000111 		: log = 32'b00000000000000001001000111001000;
			12'b110001001000 		: log = 32'b00000000000000001001000111010001;
			12'b110001001001 		: log = 32'b00000000000000001001000111011011;
			12'b110001001010 		: log = 32'b00000000000000001001000111100100;
			12'b110001001011 		: log = 32'b00000000000000001001000111101101;
			12'b110001001100 		: log = 32'b00000000000000001001000111110110;
			12'b110001001101 		: log = 32'b00000000000000001001000111111111;
			12'b110001001110 		: log = 32'b00000000000000001001001000001000;
			12'b110001001111 		: log = 32'b00000000000000001001001000010001;
			12'b110001010000 		: log = 32'b00000000000000001001001000011010;
			12'b110001010001 		: log = 32'b00000000000000001001001000100011;
			12'b110001010010 		: log = 32'b00000000000000001001001000101100;
			12'b110001010011 		: log = 32'b00000000000000001001001000110101;
			12'b110001010100 		: log = 32'b00000000000000001001001000111110;
			12'b110001010101 		: log = 32'b00000000000000001001001001000111;
			12'b110001010110 		: log = 32'b00000000000000001001001001010000;
			12'b110001010111 		: log = 32'b00000000000000001001001001011001;
			12'b110001011000 		: log = 32'b00000000000000001001001001100010;
			12'b110001011001 		: log = 32'b00000000000000001001001001101011;
			12'b110001011010 		: log = 32'b00000000000000001001001001110100;
			12'b110001011011 		: log = 32'b00000000000000001001001001111101;
			12'b110001011100 		: log = 32'b00000000000000001001001010000110;
			12'b110001011101 		: log = 32'b00000000000000001001001010001111;
			12'b110001011110 		: log = 32'b00000000000000001001001010011000;
			12'b110001011111 		: log = 32'b00000000000000001001001010100001;
			12'b110001100000 		: log = 32'b00000000000000001001001010101010;
			12'b110001100001 		: log = 32'b00000000000000001001001010110011;
			12'b110001100010 		: log = 32'b00000000000000001001001010111100;
			12'b110001100011 		: log = 32'b00000000000000001001001011000101;
			12'b110001100100 		: log = 32'b00000000000000001001001011001110;
			12'b110001100101 		: log = 32'b00000000000000001001001011010111;
			12'b110001100110 		: log = 32'b00000000000000001001001011100000;
			12'b110001100111 		: log = 32'b00000000000000001001001011101001;
			12'b110001101000 		: log = 32'b00000000000000001001001011110011;
			12'b110001101001 		: log = 32'b00000000000000001001001011111100;
			12'b110001101010 		: log = 32'b00000000000000001001001100000101;
			12'b110001101011 		: log = 32'b00000000000000001001001100001110;
			12'b110001101100 		: log = 32'b00000000000000001001001100010111;
			12'b110001101101 		: log = 32'b00000000000000001001001100100000;
			12'b110001101110 		: log = 32'b00000000000000001001001100101001;
			12'b110001101111 		: log = 32'b00000000000000001001001100110010;
			12'b110001110000 		: log = 32'b00000000000000001001001100111011;
			12'b110001110001 		: log = 32'b00000000000000001001001101000100;
			12'b110001110010 		: log = 32'b00000000000000001001001101001101;
			12'b110001110011 		: log = 32'b00000000000000001001001101010110;
			12'b110001110100 		: log = 32'b00000000000000001001001101011111;
			12'b110001110101 		: log = 32'b00000000000000001001001101101000;
			12'b110001110110 		: log = 32'b00000000000000001001001101110001;
			12'b110001110111 		: log = 32'b00000000000000001001001101111010;
			12'b110001111000 		: log = 32'b00000000000000001001001110000011;
			12'b110001111001 		: log = 32'b00000000000000001001001110001100;
			12'b110001111010 		: log = 32'b00000000000000001001001110010101;
			12'b110001111011 		: log = 32'b00000000000000001001001110011110;
			12'b110001111100 		: log = 32'b00000000000000001001001110100111;
			12'b110001111101 		: log = 32'b00000000000000001001001110101111;
			12'b110001111110 		: log = 32'b00000000000000001001001110111000;
			12'b110001111111 		: log = 32'b00000000000000001001001111000001;
			12'b110010000000 		: log = 32'b00000000000000001001001111001010;
			12'b110010000001 		: log = 32'b00000000000000001001001111010011;
			12'b110010000010 		: log = 32'b00000000000000001001001111011100;
			12'b110010000011 		: log = 32'b00000000000000001001001111100101;
			12'b110010000100 		: log = 32'b00000000000000001001001111101110;
			12'b110010000101 		: log = 32'b00000000000000001001001111110111;
			12'b110010000110 		: log = 32'b00000000000000001001010000000000;
			12'b110010000111 		: log = 32'b00000000000000001001010000001001;
			12'b110010001000 		: log = 32'b00000000000000001001010000010010;
			12'b110010001001 		: log = 32'b00000000000000001001010000011011;
			12'b110010001010 		: log = 32'b00000000000000001001010000100100;
			12'b110010001011 		: log = 32'b00000000000000001001010000101101;
			12'b110010001100 		: log = 32'b00000000000000001001010000110110;
			12'b110010001101 		: log = 32'b00000000000000001001010000111111;
			12'b110010001110 		: log = 32'b00000000000000001001010001001000;
			12'b110010001111 		: log = 32'b00000000000000001001010001010001;
			12'b110010010000 		: log = 32'b00000000000000001001010001011010;
			12'b110010010001 		: log = 32'b00000000000000001001010001100011;
			12'b110010010010 		: log = 32'b00000000000000001001010001101100;
			12'b110010010011 		: log = 32'b00000000000000001001010001110101;
			12'b110010010100 		: log = 32'b00000000000000001001010001111110;
			12'b110010010101 		: log = 32'b00000000000000001001010010000111;
			12'b110010010110 		: log = 32'b00000000000000001001010010010000;
			12'b110010010111 		: log = 32'b00000000000000001001010010011001;
			12'b110010011000 		: log = 32'b00000000000000001001010010100010;
			12'b110010011001 		: log = 32'b00000000000000001001010010101011;
			12'b110010011010 		: log = 32'b00000000000000001001010010110100;
			12'b110010011011 		: log = 32'b00000000000000001001010010111101;
			12'b110010011100 		: log = 32'b00000000000000001001010011000101;
			12'b110010011101 		: log = 32'b00000000000000001001010011001110;
			12'b110010011110 		: log = 32'b00000000000000001001010011010111;
			12'b110010011111 		: log = 32'b00000000000000001001010011100000;
			12'b110010100000 		: log = 32'b00000000000000001001010011101001;
			12'b110010100001 		: log = 32'b00000000000000001001010011110010;
			12'b110010100010 		: log = 32'b00000000000000001001010011111011;
			12'b110010100011 		: log = 32'b00000000000000001001010100000100;
			12'b110010100100 		: log = 32'b00000000000000001001010100001101;
			12'b110010100101 		: log = 32'b00000000000000001001010100010110;
			12'b110010100110 		: log = 32'b00000000000000001001010100011111;
			12'b110010100111 		: log = 32'b00000000000000001001010100101000;
			12'b110010101000 		: log = 32'b00000000000000001001010100110001;
			12'b110010101001 		: log = 32'b00000000000000001001010100111010;
			12'b110010101010 		: log = 32'b00000000000000001001010101000011;
			12'b110010101011 		: log = 32'b00000000000000001001010101001100;
			12'b110010101100 		: log = 32'b00000000000000001001010101010100;
			12'b110010101101 		: log = 32'b00000000000000001001010101011101;
			12'b110010101110 		: log = 32'b00000000000000001001010101100110;
			12'b110010101111 		: log = 32'b00000000000000001001010101101111;
			12'b110010110000 		: log = 32'b00000000000000001001010101111000;
			12'b110010110001 		: log = 32'b00000000000000001001010110000001;
			12'b110010110010 		: log = 32'b00000000000000001001010110001010;
			12'b110010110011 		: log = 32'b00000000000000001001010110010011;
			12'b110010110100 		: log = 32'b00000000000000001001010110011100;
			12'b110010110101 		: log = 32'b00000000000000001001010110100101;
			12'b110010110110 		: log = 32'b00000000000000001001010110101110;
			12'b110010110111 		: log = 32'b00000000000000001001010110110111;
			12'b110010111000 		: log = 32'b00000000000000001001010111000000;
			12'b110010111001 		: log = 32'b00000000000000001001010111001000;
			12'b110010111010 		: log = 32'b00000000000000001001010111010001;
			12'b110010111011 		: log = 32'b00000000000000001001010111011010;
			12'b110010111100 		: log = 32'b00000000000000001001010111100011;
			12'b110010111101 		: log = 32'b00000000000000001001010111101100;
			12'b110010111110 		: log = 32'b00000000000000001001010111110101;
			12'b110010111111 		: log = 32'b00000000000000001001010111111110;
			12'b110011000000 		: log = 32'b00000000000000001001011000000111;
			12'b110011000001 		: log = 32'b00000000000000001001011000010000;
			12'b110011000010 		: log = 32'b00000000000000001001011000011001;
			12'b110011000011 		: log = 32'b00000000000000001001011000100010;
			12'b110011000100 		: log = 32'b00000000000000001001011000101010;
			12'b110011000101 		: log = 32'b00000000000000001001011000110011;
			12'b110011000110 		: log = 32'b00000000000000001001011000111100;
			12'b110011000111 		: log = 32'b00000000000000001001011001000101;
			12'b110011001000 		: log = 32'b00000000000000001001011001001110;
			12'b110011001001 		: log = 32'b00000000000000001001011001010111;
			12'b110011001010 		: log = 32'b00000000000000001001011001100000;
			12'b110011001011 		: log = 32'b00000000000000001001011001101001;
			12'b110011001100 		: log = 32'b00000000000000001001011001110010;
			12'b110011001101 		: log = 32'b00000000000000001001011001111010;
			12'b110011001110 		: log = 32'b00000000000000001001011010000011;
			12'b110011001111 		: log = 32'b00000000000000001001011010001100;
			12'b110011010000 		: log = 32'b00000000000000001001011010010101;
			12'b110011010001 		: log = 32'b00000000000000001001011010011110;
			12'b110011010010 		: log = 32'b00000000000000001001011010100111;
			12'b110011010011 		: log = 32'b00000000000000001001011010110000;
			12'b110011010100 		: log = 32'b00000000000000001001011010111001;
			12'b110011010101 		: log = 32'b00000000000000001001011011000010;
			12'b110011010110 		: log = 32'b00000000000000001001011011001010;
			12'b110011010111 		: log = 32'b00000000000000001001011011010011;
			12'b110011011000 		: log = 32'b00000000000000001001011011011100;
			12'b110011011001 		: log = 32'b00000000000000001001011011100101;
			12'b110011011010 		: log = 32'b00000000000000001001011011101110;
			12'b110011011011 		: log = 32'b00000000000000001001011011110111;
			12'b110011011100 		: log = 32'b00000000000000001001011100000000;
			12'b110011011101 		: log = 32'b00000000000000001001011100001001;
			12'b110011011110 		: log = 32'b00000000000000001001011100010001;
			12'b110011011111 		: log = 32'b00000000000000001001011100011010;
			12'b110011100000 		: log = 32'b00000000000000001001011100100011;
			12'b110011100001 		: log = 32'b00000000000000001001011100101100;
			12'b110011100010 		: log = 32'b00000000000000001001011100110101;
			12'b110011100011 		: log = 32'b00000000000000001001011100111110;
			12'b110011100100 		: log = 32'b00000000000000001001011101000111;
			12'b110011100101 		: log = 32'b00000000000000001001011101001111;
			12'b110011100110 		: log = 32'b00000000000000001001011101011000;
			12'b110011100111 		: log = 32'b00000000000000001001011101100001;
			12'b110011101000 		: log = 32'b00000000000000001001011101101010;
			12'b110011101001 		: log = 32'b00000000000000001001011101110011;
			12'b110011101010 		: log = 32'b00000000000000001001011101111100;
			12'b110011101011 		: log = 32'b00000000000000001001011110000101;
			12'b110011101100 		: log = 32'b00000000000000001001011110001101;
			12'b110011101101 		: log = 32'b00000000000000001001011110010110;
			12'b110011101110 		: log = 32'b00000000000000001001011110011111;
			12'b110011101111 		: log = 32'b00000000000000001001011110101000;
			12'b110011110000 		: log = 32'b00000000000000001001011110110001;
			12'b110011110001 		: log = 32'b00000000000000001001011110111010;
			12'b110011110010 		: log = 32'b00000000000000001001011111000011;
			12'b110011110011 		: log = 32'b00000000000000001001011111001011;
			12'b110011110100 		: log = 32'b00000000000000001001011111010100;
			12'b110011110101 		: log = 32'b00000000000000001001011111011101;
			12'b110011110110 		: log = 32'b00000000000000001001011111100110;
			12'b110011110111 		: log = 32'b00000000000000001001011111101111;
			12'b110011111000 		: log = 32'b00000000000000001001011111111000;
			12'b110011111001 		: log = 32'b00000000000000001001100000000000;
			12'b110011111010 		: log = 32'b00000000000000001001100000001001;
			12'b110011111011 		: log = 32'b00000000000000001001100000010010;
			12'b110011111100 		: log = 32'b00000000000000001001100000011011;
			12'b110011111101 		: log = 32'b00000000000000001001100000100100;
			12'b110011111110 		: log = 32'b00000000000000001001100000101101;
			12'b110011111111 		: log = 32'b00000000000000001001100000110101;
			12'b110100000000 		: log = 32'b00000000000000001001100000111110;
			12'b110100000001 		: log = 32'b00000000000000001001100001000111;
			12'b110100000010 		: log = 32'b00000000000000001001100001010000;
			12'b110100000011 		: log = 32'b00000000000000001001100001011001;
			12'b110100000100 		: log = 32'b00000000000000001001100001100010;
			12'b110100000101 		: log = 32'b00000000000000001001100001101010;
			12'b110100000110 		: log = 32'b00000000000000001001100001110011;
			12'b110100000111 		: log = 32'b00000000000000001001100001111100;
			12'b110100001000 		: log = 32'b00000000000000001001100010000101;
			12'b110100001001 		: log = 32'b00000000000000001001100010001110;
			12'b110100001010 		: log = 32'b00000000000000001001100010010110;
			12'b110100001011 		: log = 32'b00000000000000001001100010011111;
			12'b110100001100 		: log = 32'b00000000000000001001100010101000;
			12'b110100001101 		: log = 32'b00000000000000001001100010110001;
			12'b110100001110 		: log = 32'b00000000000000001001100010111010;
			12'b110100001111 		: log = 32'b00000000000000001001100011000011;
			12'b110100010000 		: log = 32'b00000000000000001001100011001011;
			12'b110100010001 		: log = 32'b00000000000000001001100011010100;
			12'b110100010010 		: log = 32'b00000000000000001001100011011101;
			12'b110100010011 		: log = 32'b00000000000000001001100011100110;
			12'b110100010100 		: log = 32'b00000000000000001001100011101111;
			12'b110100010101 		: log = 32'b00000000000000001001100011110111;
			12'b110100010110 		: log = 32'b00000000000000001001100100000000;
			12'b110100010111 		: log = 32'b00000000000000001001100100001001;
			12'b110100011000 		: log = 32'b00000000000000001001100100010010;
			12'b110100011001 		: log = 32'b00000000000000001001100100011011;
			12'b110100011010 		: log = 32'b00000000000000001001100100100011;
			12'b110100011011 		: log = 32'b00000000000000001001100100101100;
			12'b110100011100 		: log = 32'b00000000000000001001100100110101;
			12'b110100011101 		: log = 32'b00000000000000001001100100111110;
			12'b110100011110 		: log = 32'b00000000000000001001100101000111;
			12'b110100011111 		: log = 32'b00000000000000001001100101001111;
			12'b110100100000 		: log = 32'b00000000000000001001100101011000;
			12'b110100100001 		: log = 32'b00000000000000001001100101100001;
			12'b110100100010 		: log = 32'b00000000000000001001100101101010;
			12'b110100100011 		: log = 32'b00000000000000001001100101110010;
			12'b110100100100 		: log = 32'b00000000000000001001100101111011;
			12'b110100100101 		: log = 32'b00000000000000001001100110000100;
			12'b110100100110 		: log = 32'b00000000000000001001100110001101;
			12'b110100100111 		: log = 32'b00000000000000001001100110010110;
			12'b110100101000 		: log = 32'b00000000000000001001100110011110;
			12'b110100101001 		: log = 32'b00000000000000001001100110100111;
			12'b110100101010 		: log = 32'b00000000000000001001100110110000;
			12'b110100101011 		: log = 32'b00000000000000001001100110111001;
			12'b110100101100 		: log = 32'b00000000000000001001100111000001;
			12'b110100101101 		: log = 32'b00000000000000001001100111001010;
			12'b110100101110 		: log = 32'b00000000000000001001100111010011;
			12'b110100101111 		: log = 32'b00000000000000001001100111011100;
			12'b110100110000 		: log = 32'b00000000000000001001100111100101;
			12'b110100110001 		: log = 32'b00000000000000001001100111101101;
			12'b110100110010 		: log = 32'b00000000000000001001100111110110;
			12'b110100110011 		: log = 32'b00000000000000001001100111111111;
			12'b110100110100 		: log = 32'b00000000000000001001101000001000;
			12'b110100110101 		: log = 32'b00000000000000001001101000010000;
			12'b110100110110 		: log = 32'b00000000000000001001101000011001;
			12'b110100110111 		: log = 32'b00000000000000001001101000100010;
			12'b110100111000 		: log = 32'b00000000000000001001101000101011;
			12'b110100111001 		: log = 32'b00000000000000001001101000110011;
			12'b110100111010 		: log = 32'b00000000000000001001101000111100;
			12'b110100111011 		: log = 32'b00000000000000001001101001000101;
			12'b110100111100 		: log = 32'b00000000000000001001101001001110;
			12'b110100111101 		: log = 32'b00000000000000001001101001010111;
			12'b110100111110 		: log = 32'b00000000000000001001101001011111;
			12'b110100111111 		: log = 32'b00000000000000001001101001101000;
			12'b110101000000 		: log = 32'b00000000000000001001101001110001;
			12'b110101000001 		: log = 32'b00000000000000001001101001111010;
			12'b110101000010 		: log = 32'b00000000000000001001101010000010;
			12'b110101000011 		: log = 32'b00000000000000001001101010001011;
			12'b110101000100 		: log = 32'b00000000000000001001101010010100;
			12'b110101000101 		: log = 32'b00000000000000001001101010011101;
			12'b110101000110 		: log = 32'b00000000000000001001101010100101;
			12'b110101000111 		: log = 32'b00000000000000001001101010101110;
			12'b110101001000 		: log = 32'b00000000000000001001101010110111;
			12'b110101001001 		: log = 32'b00000000000000001001101010111111;
			12'b110101001010 		: log = 32'b00000000000000001001101011001000;
			12'b110101001011 		: log = 32'b00000000000000001001101011010001;
			12'b110101001100 		: log = 32'b00000000000000001001101011011010;
			12'b110101001101 		: log = 32'b00000000000000001001101011100010;
			12'b110101001110 		: log = 32'b00000000000000001001101011101011;
			12'b110101001111 		: log = 32'b00000000000000001001101011110100;
			12'b110101010000 		: log = 32'b00000000000000001001101011111101;
			12'b110101010001 		: log = 32'b00000000000000001001101100000101;
			12'b110101010010 		: log = 32'b00000000000000001001101100001110;
			12'b110101010011 		: log = 32'b00000000000000001001101100010111;
			12'b110101010100 		: log = 32'b00000000000000001001101100100000;
			12'b110101010101 		: log = 32'b00000000000000001001101100101000;
			12'b110101010110 		: log = 32'b00000000000000001001101100110001;
			12'b110101010111 		: log = 32'b00000000000000001001101100111010;
			12'b110101011000 		: log = 32'b00000000000000001001101101000010;
			12'b110101011001 		: log = 32'b00000000000000001001101101001011;
			12'b110101011010 		: log = 32'b00000000000000001001101101010100;
			12'b110101011011 		: log = 32'b00000000000000001001101101011101;
			12'b110101011100 		: log = 32'b00000000000000001001101101100101;
			12'b110101011101 		: log = 32'b00000000000000001001101101101110;
			12'b110101011110 		: log = 32'b00000000000000001001101101110111;
			12'b110101011111 		: log = 32'b00000000000000001001101110000000;
			12'b110101100000 		: log = 32'b00000000000000001001101110001000;
			12'b110101100001 		: log = 32'b00000000000000001001101110010001;
			12'b110101100010 		: log = 32'b00000000000000001001101110011010;
			12'b110101100011 		: log = 32'b00000000000000001001101110100010;
			12'b110101100100 		: log = 32'b00000000000000001001101110101011;
			12'b110101100101 		: log = 32'b00000000000000001001101110110100;
			12'b110101100110 		: log = 32'b00000000000000001001101110111101;
			12'b110101100111 		: log = 32'b00000000000000001001101111000101;
			12'b110101101000 		: log = 32'b00000000000000001001101111001110;
			12'b110101101001 		: log = 32'b00000000000000001001101111010111;
			12'b110101101010 		: log = 32'b00000000000000001001101111011111;
			12'b110101101011 		: log = 32'b00000000000000001001101111101000;
			12'b110101101100 		: log = 32'b00000000000000001001101111110001;
			12'b110101101101 		: log = 32'b00000000000000001001101111111001;
			12'b110101101110 		: log = 32'b00000000000000001001110000000010;
			12'b110101101111 		: log = 32'b00000000000000001001110000001011;
			12'b110101110000 		: log = 32'b00000000000000001001110000010100;
			12'b110101110001 		: log = 32'b00000000000000001001110000011100;
			12'b110101110010 		: log = 32'b00000000000000001001110000100101;
			12'b110101110011 		: log = 32'b00000000000000001001110000101110;
			12'b110101110100 		: log = 32'b00000000000000001001110000110110;
			12'b110101110101 		: log = 32'b00000000000000001001110000111111;
			12'b110101110110 		: log = 32'b00000000000000001001110001001000;
			12'b110101110111 		: log = 32'b00000000000000001001110001010000;
			12'b110101111000 		: log = 32'b00000000000000001001110001011001;
			12'b110101111001 		: log = 32'b00000000000000001001110001100010;
			12'b110101111010 		: log = 32'b00000000000000001001110001101010;
			12'b110101111011 		: log = 32'b00000000000000001001110001110011;
			12'b110101111100 		: log = 32'b00000000000000001001110001111100;
			12'b110101111101 		: log = 32'b00000000000000001001110010000100;
			12'b110101111110 		: log = 32'b00000000000000001001110010001101;
			12'b110101111111 		: log = 32'b00000000000000001001110010010110;
			12'b110110000000 		: log = 32'b00000000000000001001110010011111;
			12'b110110000001 		: log = 32'b00000000000000001001110010100111;
			12'b110110000010 		: log = 32'b00000000000000001001110010110000;
			12'b110110000011 		: log = 32'b00000000000000001001110010111001;
			12'b110110000100 		: log = 32'b00000000000000001001110011000001;
			12'b110110000101 		: log = 32'b00000000000000001001110011001010;
			12'b110110000110 		: log = 32'b00000000000000001001110011010011;
			12'b110110000111 		: log = 32'b00000000000000001001110011011011;
			12'b110110001000 		: log = 32'b00000000000000001001110011100100;
			12'b110110001001 		: log = 32'b00000000000000001001110011101101;
			12'b110110001010 		: log = 32'b00000000000000001001110011110101;
			12'b110110001011 		: log = 32'b00000000000000001001110011111110;
			12'b110110001100 		: log = 32'b00000000000000001001110100000111;
			12'b110110001101 		: log = 32'b00000000000000001001110100001111;
			12'b110110001110 		: log = 32'b00000000000000001001110100011000;
			12'b110110001111 		: log = 32'b00000000000000001001110100100001;
			12'b110110010000 		: log = 32'b00000000000000001001110100101001;
			12'b110110010001 		: log = 32'b00000000000000001001110100110010;
			12'b110110010010 		: log = 32'b00000000000000001001110100111011;
			12'b110110010011 		: log = 32'b00000000000000001001110101000011;
			12'b110110010100 		: log = 32'b00000000000000001001110101001100;
			12'b110110010101 		: log = 32'b00000000000000001001110101010101;
			12'b110110010110 		: log = 32'b00000000000000001001110101011101;
			12'b110110010111 		: log = 32'b00000000000000001001110101100110;
			12'b110110011000 		: log = 32'b00000000000000001001110101101110;
			12'b110110011001 		: log = 32'b00000000000000001001110101110111;
			12'b110110011010 		: log = 32'b00000000000000001001110110000000;
			12'b110110011011 		: log = 32'b00000000000000001001110110001000;
			12'b110110011100 		: log = 32'b00000000000000001001110110010001;
			12'b110110011101 		: log = 32'b00000000000000001001110110011010;
			12'b110110011110 		: log = 32'b00000000000000001001110110100010;
			12'b110110011111 		: log = 32'b00000000000000001001110110101011;
			12'b110110100000 		: log = 32'b00000000000000001001110110110100;
			12'b110110100001 		: log = 32'b00000000000000001001110110111100;
			12'b110110100010 		: log = 32'b00000000000000001001110111000101;
			12'b110110100011 		: log = 32'b00000000000000001001110111001110;
			12'b110110100100 		: log = 32'b00000000000000001001110111010110;
			12'b110110100101 		: log = 32'b00000000000000001001110111011111;
			12'b110110100110 		: log = 32'b00000000000000001001110111100111;
			12'b110110100111 		: log = 32'b00000000000000001001110111110000;
			12'b110110101000 		: log = 32'b00000000000000001001110111111001;
			12'b110110101001 		: log = 32'b00000000000000001001111000000001;
			12'b110110101010 		: log = 32'b00000000000000001001111000001010;
			12'b110110101011 		: log = 32'b00000000000000001001111000010011;
			12'b110110101100 		: log = 32'b00000000000000001001111000011011;
			12'b110110101101 		: log = 32'b00000000000000001001111000100100;
			12'b110110101110 		: log = 32'b00000000000000001001111000101101;
			12'b110110101111 		: log = 32'b00000000000000001001111000110101;
			12'b110110110000 		: log = 32'b00000000000000001001111000111110;
			12'b110110110001 		: log = 32'b00000000000000001001111001000110;
			12'b110110110010 		: log = 32'b00000000000000001001111001001111;
			12'b110110110011 		: log = 32'b00000000000000001001111001011000;
			12'b110110110100 		: log = 32'b00000000000000001001111001100000;
			12'b110110110101 		: log = 32'b00000000000000001001111001101001;
			12'b110110110110 		: log = 32'b00000000000000001001111001110001;
			12'b110110110111 		: log = 32'b00000000000000001001111001111010;
			12'b110110111000 		: log = 32'b00000000000000001001111010000011;
			12'b110110111001 		: log = 32'b00000000000000001001111010001011;
			12'b110110111010 		: log = 32'b00000000000000001001111010010100;
			12'b110110111011 		: log = 32'b00000000000000001001111010011101;
			12'b110110111100 		: log = 32'b00000000000000001001111010100101;
			12'b110110111101 		: log = 32'b00000000000000001001111010101110;
			12'b110110111110 		: log = 32'b00000000000000001001111010110110;
			12'b110110111111 		: log = 32'b00000000000000001001111010111111;
			12'b110111000000 		: log = 32'b00000000000000001001111011001000;
			12'b110111000001 		: log = 32'b00000000000000001001111011010000;
			12'b110111000010 		: log = 32'b00000000000000001001111011011001;
			12'b110111000011 		: log = 32'b00000000000000001001111011100001;
			12'b110111000100 		: log = 32'b00000000000000001001111011101010;
			12'b110111000101 		: log = 32'b00000000000000001001111011110011;
			12'b110111000110 		: log = 32'b00000000000000001001111011111011;
			12'b110111000111 		: log = 32'b00000000000000001001111100000100;
			12'b110111001000 		: log = 32'b00000000000000001001111100001100;
			12'b110111001001 		: log = 32'b00000000000000001001111100010101;
			12'b110111001010 		: log = 32'b00000000000000001001111100011110;
			12'b110111001011 		: log = 32'b00000000000000001001111100100110;
			12'b110111001100 		: log = 32'b00000000000000001001111100101111;
			12'b110111001101 		: log = 32'b00000000000000001001111100110111;
			12'b110111001110 		: log = 32'b00000000000000001001111101000000;
			12'b110111001111 		: log = 32'b00000000000000001001111101001001;
			12'b110111010000 		: log = 32'b00000000000000001001111101010001;
			12'b110111010001 		: log = 32'b00000000000000001001111101011010;
			12'b110111010010 		: log = 32'b00000000000000001001111101100010;
			12'b110111010011 		: log = 32'b00000000000000001001111101101011;
			12'b110111010100 		: log = 32'b00000000000000001001111101110011;
			12'b110111010101 		: log = 32'b00000000000000001001111101111100;
			12'b110111010110 		: log = 32'b00000000000000001001111110000101;
			12'b110111010111 		: log = 32'b00000000000000001001111110001101;
			12'b110111011000 		: log = 32'b00000000000000001001111110010110;
			12'b110111011001 		: log = 32'b00000000000000001001111110011110;
			12'b110111011010 		: log = 32'b00000000000000001001111110100111;
			12'b110111011011 		: log = 32'b00000000000000001001111110110000;
			12'b110111011100 		: log = 32'b00000000000000001001111110111000;
			12'b110111011101 		: log = 32'b00000000000000001001111111000001;
			12'b110111011110 		: log = 32'b00000000000000001001111111001001;
			12'b110111011111 		: log = 32'b00000000000000001001111111010010;
			12'b110111100000 		: log = 32'b00000000000000001001111111011010;
			12'b110111100001 		: log = 32'b00000000000000001001111111100011;
			12'b110111100010 		: log = 32'b00000000000000001001111111101011;
			12'b110111100011 		: log = 32'b00000000000000001001111111110100;
			12'b110111100100 		: log = 32'b00000000000000001001111111111101;
			12'b110111100101 		: log = 32'b00000000000000001010000000000101;
			12'b110111100110 		: log = 32'b00000000000000001010000000001110;
			12'b110111100111 		: log = 32'b00000000000000001010000000010110;
			12'b110111101000 		: log = 32'b00000000000000001010000000011111;
			12'b110111101001 		: log = 32'b00000000000000001010000000100111;
			12'b110111101010 		: log = 32'b00000000000000001010000000110000;
			12'b110111101011 		: log = 32'b00000000000000001010000000111001;
			12'b110111101100 		: log = 32'b00000000000000001010000001000001;
			12'b110111101101 		: log = 32'b00000000000000001010000001001010;
			12'b110111101110 		: log = 32'b00000000000000001010000001010010;
			12'b110111101111 		: log = 32'b00000000000000001010000001011011;
			12'b110111110000 		: log = 32'b00000000000000001010000001100011;
			12'b110111110001 		: log = 32'b00000000000000001010000001101100;
			12'b110111110010 		: log = 32'b00000000000000001010000001110100;
			12'b110111110011 		: log = 32'b00000000000000001010000001111101;
			12'b110111110100 		: log = 32'b00000000000000001010000010000110;
			12'b110111110101 		: log = 32'b00000000000000001010000010001110;
			12'b110111110110 		: log = 32'b00000000000000001010000010010111;
			12'b110111110111 		: log = 32'b00000000000000001010000010011111;
			12'b110111111000 		: log = 32'b00000000000000001010000010101000;
			12'b110111111001 		: log = 32'b00000000000000001010000010110000;
			12'b110111111010 		: log = 32'b00000000000000001010000010111001;
			12'b110111111011 		: log = 32'b00000000000000001010000011000001;
			12'b110111111100 		: log = 32'b00000000000000001010000011001010;
			12'b110111111101 		: log = 32'b00000000000000001010000011010010;
			12'b110111111110 		: log = 32'b00000000000000001010000011011011;
			12'b110111111111 		: log = 32'b00000000000000001010000011100011;
			12'b111000000000 		: log = 32'b00000000000000001010000011101100;
			12'b111000000001 		: log = 32'b00000000000000001010000011110101;
			12'b111000000010 		: log = 32'b00000000000000001010000011111101;
			12'b111000000011 		: log = 32'b00000000000000001010000100000110;
			12'b111000000100 		: log = 32'b00000000000000001010000100001110;
			12'b111000000101 		: log = 32'b00000000000000001010000100010111;
			12'b111000000110 		: log = 32'b00000000000000001010000100011111;
			12'b111000000111 		: log = 32'b00000000000000001010000100101000;
			12'b111000001000 		: log = 32'b00000000000000001010000100110000;
			12'b111000001001 		: log = 32'b00000000000000001010000100111001;
			12'b111000001010 		: log = 32'b00000000000000001010000101000001;
			12'b111000001011 		: log = 32'b00000000000000001010000101001010;
			12'b111000001100 		: log = 32'b00000000000000001010000101010010;
			12'b111000001101 		: log = 32'b00000000000000001010000101011011;
			12'b111000001110 		: log = 32'b00000000000000001010000101100011;
			12'b111000001111 		: log = 32'b00000000000000001010000101101100;
			12'b111000010000 		: log = 32'b00000000000000001010000101110100;
			12'b111000010001 		: log = 32'b00000000000000001010000101111101;
			12'b111000010010 		: log = 32'b00000000000000001010000110000101;
			12'b111000010011 		: log = 32'b00000000000000001010000110001110;
			12'b111000010100 		: log = 32'b00000000000000001010000110010110;
			12'b111000010101 		: log = 32'b00000000000000001010000110011111;
			12'b111000010110 		: log = 32'b00000000000000001010000110100111;
			12'b111000010111 		: log = 32'b00000000000000001010000110110000;
			12'b111000011000 		: log = 32'b00000000000000001010000110111000;
			12'b111000011001 		: log = 32'b00000000000000001010000111000001;
			12'b111000011010 		: log = 32'b00000000000000001010000111001001;
			12'b111000011011 		: log = 32'b00000000000000001010000111010010;
			12'b111000011100 		: log = 32'b00000000000000001010000111011010;
			12'b111000011101 		: log = 32'b00000000000000001010000111100011;
			12'b111000011110 		: log = 32'b00000000000000001010000111101011;
			12'b111000011111 		: log = 32'b00000000000000001010000111110100;
			12'b111000100000 		: log = 32'b00000000000000001010000111111100;
			12'b111000100001 		: log = 32'b00000000000000001010001000000101;
			12'b111000100010 		: log = 32'b00000000000000001010001000001101;
			12'b111000100011 		: log = 32'b00000000000000001010001000010110;
			12'b111000100100 		: log = 32'b00000000000000001010001000011110;
			12'b111000100101 		: log = 32'b00000000000000001010001000100111;
			12'b111000100110 		: log = 32'b00000000000000001010001000101111;
			12'b111000100111 		: log = 32'b00000000000000001010001000111000;
			12'b111000101000 		: log = 32'b00000000000000001010001001000000;
			12'b111000101001 		: log = 32'b00000000000000001010001001001001;
			12'b111000101010 		: log = 32'b00000000000000001010001001010001;
			12'b111000101011 		: log = 32'b00000000000000001010001001011010;
			12'b111000101100 		: log = 32'b00000000000000001010001001100010;
			12'b111000101101 		: log = 32'b00000000000000001010001001101011;
			12'b111000101110 		: log = 32'b00000000000000001010001001110011;
			12'b111000101111 		: log = 32'b00000000000000001010001001111100;
			12'b111000110000 		: log = 32'b00000000000000001010001010000100;
			12'b111000110001 		: log = 32'b00000000000000001010001010001101;
			12'b111000110010 		: log = 32'b00000000000000001010001010010101;
			12'b111000110011 		: log = 32'b00000000000000001010001010011110;
			12'b111000110100 		: log = 32'b00000000000000001010001010100110;
			12'b111000110101 		: log = 32'b00000000000000001010001010101111;
			12'b111000110110 		: log = 32'b00000000000000001010001010110111;
			12'b111000110111 		: log = 32'b00000000000000001010001011000000;
			12'b111000111000 		: log = 32'b00000000000000001010001011001000;
			12'b111000111001 		: log = 32'b00000000000000001010001011010001;
			12'b111000111010 		: log = 32'b00000000000000001010001011011001;
			12'b111000111011 		: log = 32'b00000000000000001010001011100010;
			12'b111000111100 		: log = 32'b00000000000000001010001011101010;
			12'b111000111101 		: log = 32'b00000000000000001010001011110010;
			12'b111000111110 		: log = 32'b00000000000000001010001011111011;
			12'b111000111111 		: log = 32'b00000000000000001010001100000011;
			12'b111001000000 		: log = 32'b00000000000000001010001100001100;
			12'b111001000001 		: log = 32'b00000000000000001010001100010100;
			12'b111001000010 		: log = 32'b00000000000000001010001100011101;
			12'b111001000011 		: log = 32'b00000000000000001010001100100101;
			12'b111001000100 		: log = 32'b00000000000000001010001100101110;
			12'b111001000101 		: log = 32'b00000000000000001010001100110110;
			12'b111001000110 		: log = 32'b00000000000000001010001100111111;
			12'b111001000111 		: log = 32'b00000000000000001010001101000111;
			12'b111001001000 		: log = 32'b00000000000000001010001101010000;
			12'b111001001001 		: log = 32'b00000000000000001010001101011000;
			12'b111001001010 		: log = 32'b00000000000000001010001101100000;
			12'b111001001011 		: log = 32'b00000000000000001010001101101001;
			12'b111001001100 		: log = 32'b00000000000000001010001101110001;
			12'b111001001101 		: log = 32'b00000000000000001010001101111010;
			12'b111001001110 		: log = 32'b00000000000000001010001110000010;
			12'b111001001111 		: log = 32'b00000000000000001010001110001011;
			12'b111001010000 		: log = 32'b00000000000000001010001110010011;
			12'b111001010001 		: log = 32'b00000000000000001010001110011100;
			12'b111001010010 		: log = 32'b00000000000000001010001110100100;
			12'b111001010011 		: log = 32'b00000000000000001010001110101100;
			12'b111001010100 		: log = 32'b00000000000000001010001110110101;
			12'b111001010101 		: log = 32'b00000000000000001010001110111101;
			12'b111001010110 		: log = 32'b00000000000000001010001111000110;
			12'b111001010111 		: log = 32'b00000000000000001010001111001110;
			12'b111001011000 		: log = 32'b00000000000000001010001111010111;
			12'b111001011001 		: log = 32'b00000000000000001010001111011111;
			12'b111001011010 		: log = 32'b00000000000000001010001111101000;
			12'b111001011011 		: log = 32'b00000000000000001010001111110000;
			12'b111001011100 		: log = 32'b00000000000000001010001111111000;
			12'b111001011101 		: log = 32'b00000000000000001010010000000001;
			12'b111001011110 		: log = 32'b00000000000000001010010000001001;
			12'b111001011111 		: log = 32'b00000000000000001010010000010010;
			12'b111001100000 		: log = 32'b00000000000000001010010000011010;
			12'b111001100001 		: log = 32'b00000000000000001010010000100011;
			12'b111001100010 		: log = 32'b00000000000000001010010000101011;
			12'b111001100011 		: log = 32'b00000000000000001010010000110011;
			12'b111001100100 		: log = 32'b00000000000000001010010000111100;
			12'b111001100101 		: log = 32'b00000000000000001010010001000100;
			12'b111001100110 		: log = 32'b00000000000000001010010001001101;
			12'b111001100111 		: log = 32'b00000000000000001010010001010101;
			12'b111001101000 		: log = 32'b00000000000000001010010001011110;
			12'b111001101001 		: log = 32'b00000000000000001010010001100110;
			12'b111001101010 		: log = 32'b00000000000000001010010001101110;
			12'b111001101011 		: log = 32'b00000000000000001010010001110111;
			12'b111001101100 		: log = 32'b00000000000000001010010001111111;
			12'b111001101101 		: log = 32'b00000000000000001010010010001000;
			12'b111001101110 		: log = 32'b00000000000000001010010010010000;
			12'b111001101111 		: log = 32'b00000000000000001010010010011000;
			12'b111001110000 		: log = 32'b00000000000000001010010010100001;
			12'b111001110001 		: log = 32'b00000000000000001010010010101001;
			12'b111001110010 		: log = 32'b00000000000000001010010010110010;
			12'b111001110011 		: log = 32'b00000000000000001010010010111010;
			12'b111001110100 		: log = 32'b00000000000000001010010011000010;
			12'b111001110101 		: log = 32'b00000000000000001010010011001011;
			12'b111001110110 		: log = 32'b00000000000000001010010011010011;
			12'b111001110111 		: log = 32'b00000000000000001010010011011100;
			12'b111001111000 		: log = 32'b00000000000000001010010011100100;
			12'b111001111001 		: log = 32'b00000000000000001010010011101100;
			12'b111001111010 		: log = 32'b00000000000000001010010011110101;
			12'b111001111011 		: log = 32'b00000000000000001010010011111101;
			12'b111001111100 		: log = 32'b00000000000000001010010100000110;
			12'b111001111101 		: log = 32'b00000000000000001010010100001110;
			12'b111001111110 		: log = 32'b00000000000000001010010100010110;
			12'b111001111111 		: log = 32'b00000000000000001010010100011111;
			12'b111010000000 		: log = 32'b00000000000000001010010100100111;
			12'b111010000001 		: log = 32'b00000000000000001010010100110000;
			12'b111010000010 		: log = 32'b00000000000000001010010100111000;
			12'b111010000011 		: log = 32'b00000000000000001010010101000000;
			12'b111010000100 		: log = 32'b00000000000000001010010101001001;
			12'b111010000101 		: log = 32'b00000000000000001010010101010001;
			12'b111010000110 		: log = 32'b00000000000000001010010101011010;
			12'b111010000111 		: log = 32'b00000000000000001010010101100010;
			12'b111010001000 		: log = 32'b00000000000000001010010101101010;
			12'b111010001001 		: log = 32'b00000000000000001010010101110011;
			12'b111010001010 		: log = 32'b00000000000000001010010101111011;
			12'b111010001011 		: log = 32'b00000000000000001010010110000100;
			12'b111010001100 		: log = 32'b00000000000000001010010110001100;
			12'b111010001101 		: log = 32'b00000000000000001010010110010100;
			12'b111010001110 		: log = 32'b00000000000000001010010110011101;
			12'b111010001111 		: log = 32'b00000000000000001010010110100101;
			12'b111010010000 		: log = 32'b00000000000000001010010110101101;
			12'b111010010001 		: log = 32'b00000000000000001010010110110110;
			12'b111010010010 		: log = 32'b00000000000000001010010110111110;
			12'b111010010011 		: log = 32'b00000000000000001010010111000111;
			12'b111010010100 		: log = 32'b00000000000000001010010111001111;
			12'b111010010101 		: log = 32'b00000000000000001010010111010111;
			12'b111010010110 		: log = 32'b00000000000000001010010111100000;
			12'b111010010111 		: log = 32'b00000000000000001010010111101000;
			12'b111010011000 		: log = 32'b00000000000000001010010111110000;
			12'b111010011001 		: log = 32'b00000000000000001010010111111001;
			12'b111010011010 		: log = 32'b00000000000000001010011000000001;
			12'b111010011011 		: log = 32'b00000000000000001010011000001001;
			12'b111010011100 		: log = 32'b00000000000000001010011000010010;
			12'b111010011101 		: log = 32'b00000000000000001010011000011010;
			12'b111010011110 		: log = 32'b00000000000000001010011000100011;
			12'b111010011111 		: log = 32'b00000000000000001010011000101011;
			12'b111010100000 		: log = 32'b00000000000000001010011000110011;
			12'b111010100001 		: log = 32'b00000000000000001010011000111100;
			12'b111010100010 		: log = 32'b00000000000000001010011001000100;
			12'b111010100011 		: log = 32'b00000000000000001010011001001100;
			12'b111010100100 		: log = 32'b00000000000000001010011001010101;
			12'b111010100101 		: log = 32'b00000000000000001010011001011101;
			12'b111010100110 		: log = 32'b00000000000000001010011001100101;
			12'b111010100111 		: log = 32'b00000000000000001010011001101110;
			12'b111010101000 		: log = 32'b00000000000000001010011001110110;
			12'b111010101001 		: log = 32'b00000000000000001010011001111110;
			12'b111010101010 		: log = 32'b00000000000000001010011010000111;
			12'b111010101011 		: log = 32'b00000000000000001010011010001111;
			12'b111010101100 		: log = 32'b00000000000000001010011010011000;
			12'b111010101101 		: log = 32'b00000000000000001010011010100000;
			12'b111010101110 		: log = 32'b00000000000000001010011010101000;
			12'b111010101111 		: log = 32'b00000000000000001010011010110001;
			12'b111010110000 		: log = 32'b00000000000000001010011010111001;
			12'b111010110001 		: log = 32'b00000000000000001010011011000001;
			12'b111010110010 		: log = 32'b00000000000000001010011011001010;
			12'b111010110011 		: log = 32'b00000000000000001010011011010010;
			12'b111010110100 		: log = 32'b00000000000000001010011011011010;
			12'b111010110101 		: log = 32'b00000000000000001010011011100011;
			12'b111010110110 		: log = 32'b00000000000000001010011011101011;
			12'b111010110111 		: log = 32'b00000000000000001010011011110011;
			12'b111010111000 		: log = 32'b00000000000000001010011011111100;
			12'b111010111001 		: log = 32'b00000000000000001010011100000100;
			12'b111010111010 		: log = 32'b00000000000000001010011100001100;
			12'b111010111011 		: log = 32'b00000000000000001010011100010101;
			12'b111010111100 		: log = 32'b00000000000000001010011100011101;
			12'b111010111101 		: log = 32'b00000000000000001010011100100101;
			12'b111010111110 		: log = 32'b00000000000000001010011100101110;
			12'b111010111111 		: log = 32'b00000000000000001010011100110110;
			12'b111011000000 		: log = 32'b00000000000000001010011100111110;
			12'b111011000001 		: log = 32'b00000000000000001010011101000111;
			12'b111011000010 		: log = 32'b00000000000000001010011101001111;
			12'b111011000011 		: log = 32'b00000000000000001010011101010111;
			12'b111011000100 		: log = 32'b00000000000000001010011101100000;
			12'b111011000101 		: log = 32'b00000000000000001010011101101000;
			12'b111011000110 		: log = 32'b00000000000000001010011101110000;
			12'b111011000111 		: log = 32'b00000000000000001010011101111001;
			12'b111011001000 		: log = 32'b00000000000000001010011110000001;
			12'b111011001001 		: log = 32'b00000000000000001010011110001001;
			12'b111011001010 		: log = 32'b00000000000000001010011110010001;
			12'b111011001011 		: log = 32'b00000000000000001010011110011010;
			12'b111011001100 		: log = 32'b00000000000000001010011110100010;
			12'b111011001101 		: log = 32'b00000000000000001010011110101010;
			12'b111011001110 		: log = 32'b00000000000000001010011110110011;
			12'b111011001111 		: log = 32'b00000000000000001010011110111011;
			12'b111011010000 		: log = 32'b00000000000000001010011111000011;
			12'b111011010001 		: log = 32'b00000000000000001010011111001100;
			12'b111011010010 		: log = 32'b00000000000000001010011111010100;
			12'b111011010011 		: log = 32'b00000000000000001010011111011100;
			12'b111011010100 		: log = 32'b00000000000000001010011111100101;
			12'b111011010101 		: log = 32'b00000000000000001010011111101101;
			12'b111011010110 		: log = 32'b00000000000000001010011111110101;
			12'b111011010111 		: log = 32'b00000000000000001010011111111101;
			12'b111011011000 		: log = 32'b00000000000000001010100000000110;
			12'b111011011001 		: log = 32'b00000000000000001010100000001110;
			12'b111011011010 		: log = 32'b00000000000000001010100000010110;
			12'b111011011011 		: log = 32'b00000000000000001010100000011111;
			12'b111011011100 		: log = 32'b00000000000000001010100000100111;
			12'b111011011101 		: log = 32'b00000000000000001010100000101111;
			12'b111011011110 		: log = 32'b00000000000000001010100000111000;
			12'b111011011111 		: log = 32'b00000000000000001010100001000000;
			12'b111011100000 		: log = 32'b00000000000000001010100001001000;
			12'b111011100001 		: log = 32'b00000000000000001010100001010000;
			12'b111011100010 		: log = 32'b00000000000000001010100001011001;
			12'b111011100011 		: log = 32'b00000000000000001010100001100001;
			12'b111011100100 		: log = 32'b00000000000000001010100001101001;
			12'b111011100101 		: log = 32'b00000000000000001010100001110010;
			12'b111011100110 		: log = 32'b00000000000000001010100001111010;
			12'b111011100111 		: log = 32'b00000000000000001010100010000010;
			12'b111011101000 		: log = 32'b00000000000000001010100010001010;
			12'b111011101001 		: log = 32'b00000000000000001010100010010011;
			12'b111011101010 		: log = 32'b00000000000000001010100010011011;
			12'b111011101011 		: log = 32'b00000000000000001010100010100011;
			12'b111011101100 		: log = 32'b00000000000000001010100010101100;
			12'b111011101101 		: log = 32'b00000000000000001010100010110100;
			12'b111011101110 		: log = 32'b00000000000000001010100010111100;
			12'b111011101111 		: log = 32'b00000000000000001010100011000100;
			12'b111011110000 		: log = 32'b00000000000000001010100011001101;
			12'b111011110001 		: log = 32'b00000000000000001010100011010101;
			12'b111011110010 		: log = 32'b00000000000000001010100011011101;
			12'b111011110011 		: log = 32'b00000000000000001010100011100101;
			12'b111011110100 		: log = 32'b00000000000000001010100011101110;
			12'b111011110101 		: log = 32'b00000000000000001010100011110110;
			12'b111011110110 		: log = 32'b00000000000000001010100011111110;
			12'b111011110111 		: log = 32'b00000000000000001010100100000111;
			12'b111011111000 		: log = 32'b00000000000000001010100100001111;
			12'b111011111001 		: log = 32'b00000000000000001010100100010111;
			12'b111011111010 		: log = 32'b00000000000000001010100100011111;
			12'b111011111011 		: log = 32'b00000000000000001010100100101000;
			12'b111011111100 		: log = 32'b00000000000000001010100100110000;
			12'b111011111101 		: log = 32'b00000000000000001010100100111000;
			12'b111011111110 		: log = 32'b00000000000000001010100101000000;
			12'b111011111111 		: log = 32'b00000000000000001010100101001001;
			12'b111100000000 		: log = 32'b00000000000000001010100101010001;
			12'b111100000001 		: log = 32'b00000000000000001010100101011001;
			12'b111100000010 		: log = 32'b00000000000000001010100101100001;
			12'b111100000011 		: log = 32'b00000000000000001010100101101010;
			12'b111100000100 		: log = 32'b00000000000000001010100101110010;
			12'b111100000101 		: log = 32'b00000000000000001010100101111010;
			12'b111100000110 		: log = 32'b00000000000000001010100110000010;
			12'b111100000111 		: log = 32'b00000000000000001010100110001011;
			12'b111100001000 		: log = 32'b00000000000000001010100110010011;
			12'b111100001001 		: log = 32'b00000000000000001010100110011011;
			12'b111100001010 		: log = 32'b00000000000000001010100110100011;
			12'b111100001011 		: log = 32'b00000000000000001010100110101100;
			12'b111100001100 		: log = 32'b00000000000000001010100110110100;
			12'b111100001101 		: log = 32'b00000000000000001010100110111100;
			12'b111100001110 		: log = 32'b00000000000000001010100111000100;
			12'b111100001111 		: log = 32'b00000000000000001010100111001101;
			12'b111100010000 		: log = 32'b00000000000000001010100111010101;
			12'b111100010001 		: log = 32'b00000000000000001010100111011101;
			12'b111100010010 		: log = 32'b00000000000000001010100111100101;
			12'b111100010011 		: log = 32'b00000000000000001010100111101110;
			12'b111100010100 		: log = 32'b00000000000000001010100111110110;
			12'b111100010101 		: log = 32'b00000000000000001010100111111110;
			12'b111100010110 		: log = 32'b00000000000000001010101000000110;
			12'b111100010111 		: log = 32'b00000000000000001010101000001111;
			12'b111100011000 		: log = 32'b00000000000000001010101000010111;
			12'b111100011001 		: log = 32'b00000000000000001010101000011111;
			12'b111100011010 		: log = 32'b00000000000000001010101000100111;
			12'b111100011011 		: log = 32'b00000000000000001010101000110000;
			12'b111100011100 		: log = 32'b00000000000000001010101000111000;
			12'b111100011101 		: log = 32'b00000000000000001010101001000000;
			12'b111100011110 		: log = 32'b00000000000000001010101001001000;
			12'b111100011111 		: log = 32'b00000000000000001010101001010000;
			12'b111100100000 		: log = 32'b00000000000000001010101001011001;
			12'b111100100001 		: log = 32'b00000000000000001010101001100001;
			12'b111100100010 		: log = 32'b00000000000000001010101001101001;
			12'b111100100011 		: log = 32'b00000000000000001010101001110001;
			12'b111100100100 		: log = 32'b00000000000000001010101001111010;
			12'b111100100101 		: log = 32'b00000000000000001010101010000010;
			12'b111100100110 		: log = 32'b00000000000000001010101010001010;
			12'b111100100111 		: log = 32'b00000000000000001010101010010010;
			12'b111100101000 		: log = 32'b00000000000000001010101010011010;
			12'b111100101001 		: log = 32'b00000000000000001010101010100011;
			12'b111100101010 		: log = 32'b00000000000000001010101010101011;
			12'b111100101011 		: log = 32'b00000000000000001010101010110011;
			12'b111100101100 		: log = 32'b00000000000000001010101010111011;
			12'b111100101101 		: log = 32'b00000000000000001010101011000011;
			12'b111100101110 		: log = 32'b00000000000000001010101011001100;
			12'b111100101111 		: log = 32'b00000000000000001010101011010100;
			12'b111100110000 		: log = 32'b00000000000000001010101011011100;
			12'b111100110001 		: log = 32'b00000000000000001010101011100100;
			12'b111100110010 		: log = 32'b00000000000000001010101011101101;
			12'b111100110011 		: log = 32'b00000000000000001010101011110101;
			12'b111100110100 		: log = 32'b00000000000000001010101011111101;
			12'b111100110101 		: log = 32'b00000000000000001010101100000101;
			12'b111100110110 		: log = 32'b00000000000000001010101100001101;
			12'b111100110111 		: log = 32'b00000000000000001010101100010110;
			12'b111100111000 		: log = 32'b00000000000000001010101100011110;
			12'b111100111001 		: log = 32'b00000000000000001010101100100110;
			12'b111100111010 		: log = 32'b00000000000000001010101100101110;
			12'b111100111011 		: log = 32'b00000000000000001010101100110110;
			12'b111100111100 		: log = 32'b00000000000000001010101100111111;
			12'b111100111101 		: log = 32'b00000000000000001010101101000111;
			12'b111100111110 		: log = 32'b00000000000000001010101101001111;
			12'b111100111111 		: log = 32'b00000000000000001010101101010111;
			12'b111101000000 		: log = 32'b00000000000000001010101101011111;
			12'b111101000001 		: log = 32'b00000000000000001010101101100111;
			12'b111101000010 		: log = 32'b00000000000000001010101101110000;
			12'b111101000011 		: log = 32'b00000000000000001010101101111000;
			12'b111101000100 		: log = 32'b00000000000000001010101110000000;
			12'b111101000101 		: log = 32'b00000000000000001010101110001000;
			12'b111101000110 		: log = 32'b00000000000000001010101110010000;
			12'b111101000111 		: log = 32'b00000000000000001010101110011001;
			12'b111101001000 		: log = 32'b00000000000000001010101110100001;
			12'b111101001001 		: log = 32'b00000000000000001010101110101001;
			12'b111101001010 		: log = 32'b00000000000000001010101110110001;
			12'b111101001011 		: log = 32'b00000000000000001010101110111001;
			12'b111101001100 		: log = 32'b00000000000000001010101111000010;
			12'b111101001101 		: log = 32'b00000000000000001010101111001010;
			12'b111101001110 		: log = 32'b00000000000000001010101111010010;
			12'b111101001111 		: log = 32'b00000000000000001010101111011010;
			12'b111101010000 		: log = 32'b00000000000000001010101111100010;
			12'b111101010001 		: log = 32'b00000000000000001010101111101010;
			12'b111101010010 		: log = 32'b00000000000000001010101111110011;
			12'b111101010011 		: log = 32'b00000000000000001010101111111011;
			12'b111101010100 		: log = 32'b00000000000000001010110000000011;
			12'b111101010101 		: log = 32'b00000000000000001010110000001011;
			12'b111101010110 		: log = 32'b00000000000000001010110000010011;
			12'b111101010111 		: log = 32'b00000000000000001010110000011011;
			12'b111101011000 		: log = 32'b00000000000000001010110000100100;
			12'b111101011001 		: log = 32'b00000000000000001010110000101100;
			12'b111101011010 		: log = 32'b00000000000000001010110000110100;
			12'b111101011011 		: log = 32'b00000000000000001010110000111100;
			12'b111101011100 		: log = 32'b00000000000000001010110001000100;
			12'b111101011101 		: log = 32'b00000000000000001010110001001100;
			12'b111101011110 		: log = 32'b00000000000000001010110001010101;
			12'b111101011111 		: log = 32'b00000000000000001010110001011101;
			12'b111101100000 		: log = 32'b00000000000000001010110001100101;
			12'b111101100001 		: log = 32'b00000000000000001010110001101101;
			12'b111101100010 		: log = 32'b00000000000000001010110001110101;
			12'b111101100011 		: log = 32'b00000000000000001010110001111101;
			12'b111101100100 		: log = 32'b00000000000000001010110010000110;
			12'b111101100101 		: log = 32'b00000000000000001010110010001110;
			12'b111101100110 		: log = 32'b00000000000000001010110010010110;
			12'b111101100111 		: log = 32'b00000000000000001010110010011110;
			12'b111101101000 		: log = 32'b00000000000000001010110010100110;
			12'b111101101001 		: log = 32'b00000000000000001010110010101110;
			12'b111101101010 		: log = 32'b00000000000000001010110010110110;
			12'b111101101011 		: log = 32'b00000000000000001010110010111111;
			12'b111101101100 		: log = 32'b00000000000000001010110011000111;
			12'b111101101101 		: log = 32'b00000000000000001010110011001111;
			12'b111101101110 		: log = 32'b00000000000000001010110011010111;
			12'b111101101111 		: log = 32'b00000000000000001010110011011111;
			12'b111101110000 		: log = 32'b00000000000000001010110011100111;
			12'b111101110001 		: log = 32'b00000000000000001010110011101111;
			12'b111101110010 		: log = 32'b00000000000000001010110011111000;
			12'b111101110011 		: log = 32'b00000000000000001010110100000000;
			12'b111101110100 		: log = 32'b00000000000000001010110100001000;
			12'b111101110101 		: log = 32'b00000000000000001010110100010000;
			12'b111101110110 		: log = 32'b00000000000000001010110100011000;
			12'b111101110111 		: log = 32'b00000000000000001010110100100000;
			12'b111101111000 		: log = 32'b00000000000000001010110100101000;
			12'b111101111001 		: log = 32'b00000000000000001010110100110001;
			12'b111101111010 		: log = 32'b00000000000000001010110100111001;
			12'b111101111011 		: log = 32'b00000000000000001010110101000001;
			12'b111101111100 		: log = 32'b00000000000000001010110101001001;
			12'b111101111101 		: log = 32'b00000000000000001010110101010001;
			12'b111101111110 		: log = 32'b00000000000000001010110101011001;
			12'b111101111111 		: log = 32'b00000000000000001010110101100001;
			12'b111110000000 		: log = 32'b00000000000000001010110101101010;
			12'b111110000001 		: log = 32'b00000000000000001010110101110010;
			12'b111110000010 		: log = 32'b00000000000000001010110101111010;
			12'b111110000011 		: log = 32'b00000000000000001010110110000010;
			12'b111110000100 		: log = 32'b00000000000000001010110110001010;
			12'b111110000101 		: log = 32'b00000000000000001010110110010010;
			12'b111110000110 		: log = 32'b00000000000000001010110110011010;
			12'b111110000111 		: log = 32'b00000000000000001010110110100010;
			12'b111110001000 		: log = 32'b00000000000000001010110110101010;
			12'b111110001001 		: log = 32'b00000000000000001010110110110011;
			12'b111110001010 		: log = 32'b00000000000000001010110110111011;
			12'b111110001011 		: log = 32'b00000000000000001010110111000011;
			12'b111110001100 		: log = 32'b00000000000000001010110111001011;
			12'b111110001101 		: log = 32'b00000000000000001010110111010011;
			12'b111110001110 		: log = 32'b00000000000000001010110111011011;
			12'b111110001111 		: log = 32'b00000000000000001010110111100011;
			12'b111110010000 		: log = 32'b00000000000000001010110111101011;
			12'b111110010001 		: log = 32'b00000000000000001010110111110100;
			12'b111110010010 		: log = 32'b00000000000000001010110111111100;
			12'b111110010011 		: log = 32'b00000000000000001010111000000100;
			12'b111110010100 		: log = 32'b00000000000000001010111000001100;
			12'b111110010101 		: log = 32'b00000000000000001010111000010100;
			12'b111110010110 		: log = 32'b00000000000000001010111000011100;
			12'b111110010111 		: log = 32'b00000000000000001010111000100100;
			12'b111110011000 		: log = 32'b00000000000000001010111000101100;
			12'b111110011001 		: log = 32'b00000000000000001010111000110100;
			12'b111110011010 		: log = 32'b00000000000000001010111000111100;
			12'b111110011011 		: log = 32'b00000000000000001010111001000101;
			12'b111110011100 		: log = 32'b00000000000000001010111001001101;
			12'b111110011101 		: log = 32'b00000000000000001010111001010101;
			12'b111110011110 		: log = 32'b00000000000000001010111001011101;
			12'b111110011111 		: log = 32'b00000000000000001010111001100101;
			12'b111110100000 		: log = 32'b00000000000000001010111001101101;
			12'b111110100001 		: log = 32'b00000000000000001010111001110101;
			12'b111110100010 		: log = 32'b00000000000000001010111001111101;
			12'b111110100011 		: log = 32'b00000000000000001010111010000101;
			12'b111110100100 		: log = 32'b00000000000000001010111010001101;
			12'b111110100101 		: log = 32'b00000000000000001010111010010110;
			12'b111110100110 		: log = 32'b00000000000000001010111010011110;
			12'b111110100111 		: log = 32'b00000000000000001010111010100110;
			12'b111110101000 		: log = 32'b00000000000000001010111010101110;
			12'b111110101001 		: log = 32'b00000000000000001010111010110110;
			12'b111110101010 		: log = 32'b00000000000000001010111010111110;
			12'b111110101011 		: log = 32'b00000000000000001010111011000110;
			12'b111110101100 		: log = 32'b00000000000000001010111011001110;
			12'b111110101101 		: log = 32'b00000000000000001010111011010110;
			12'b111110101110 		: log = 32'b00000000000000001010111011011110;
			12'b111110101111 		: log = 32'b00000000000000001010111011100110;
			12'b111110110000 		: log = 32'b00000000000000001010111011101110;
			12'b111110110001 		: log = 32'b00000000000000001010111011110111;
			12'b111110110010 		: log = 32'b00000000000000001010111011111111;
			12'b111110110011 		: log = 32'b00000000000000001010111100000111;
			12'b111110110100 		: log = 32'b00000000000000001010111100001111;
			12'b111110110101 		: log = 32'b00000000000000001010111100010111;
			12'b111110110110 		: log = 32'b00000000000000001010111100011111;
			12'b111110110111 		: log = 32'b00000000000000001010111100100111;
			12'b111110111000 		: log = 32'b00000000000000001010111100101111;
			12'b111110111001 		: log = 32'b00000000000000001010111100110111;
			12'b111110111010 		: log = 32'b00000000000000001010111100111111;
			12'b111110111011 		: log = 32'b00000000000000001010111101000111;
			12'b111110111100 		: log = 32'b00000000000000001010111101001111;
			12'b111110111101 		: log = 32'b00000000000000001010111101010111;
			12'b111110111110 		: log = 32'b00000000000000001010111101011111;
			12'b111110111111 		: log = 32'b00000000000000001010111101101000;
			12'b111111000000 		: log = 32'b00000000000000001010111101110000;
			12'b111111000001 		: log = 32'b00000000000000001010111101111000;
			12'b111111000010 		: log = 32'b00000000000000001010111110000000;
			12'b111111000011 		: log = 32'b00000000000000001010111110001000;
			12'b111111000100 		: log = 32'b00000000000000001010111110010000;
			12'b111111000101 		: log = 32'b00000000000000001010111110011000;
			12'b111111000110 		: log = 32'b00000000000000001010111110100000;
			12'b111111000111 		: log = 32'b00000000000000001010111110101000;
			12'b111111001000 		: log = 32'b00000000000000001010111110110000;
			12'b111111001001 		: log = 32'b00000000000000001010111110111000;
			12'b111111001010 		: log = 32'b00000000000000001010111111000000;
			12'b111111001011 		: log = 32'b00000000000000001010111111001000;
			12'b111111001100 		: log = 32'b00000000000000001010111111010000;
			12'b111111001101 		: log = 32'b00000000000000001010111111011000;
			12'b111111001110 		: log = 32'b00000000000000001010111111100000;
			12'b111111001111 		: log = 32'b00000000000000001010111111101000;
			12'b111111010000 		: log = 32'b00000000000000001010111111110000;
			12'b111111010001 		: log = 32'b00000000000000001010111111111001;
			12'b111111010010 		: log = 32'b00000000000000001011000000000001;
			12'b111111010011 		: log = 32'b00000000000000001011000000001001;
			12'b111111010100 		: log = 32'b00000000000000001011000000010001;
			12'b111111010101 		: log = 32'b00000000000000001011000000011001;
			12'b111111010110 		: log = 32'b00000000000000001011000000100001;
			12'b111111010111 		: log = 32'b00000000000000001011000000101001;
			12'b111111011000 		: log = 32'b00000000000000001011000000110001;
			12'b111111011001 		: log = 32'b00000000000000001011000000111001;
			12'b111111011010 		: log = 32'b00000000000000001011000001000001;
			12'b111111011011 		: log = 32'b00000000000000001011000001001001;
			12'b111111011100 		: log = 32'b00000000000000001011000001010001;
			12'b111111011101 		: log = 32'b00000000000000001011000001011001;
			12'b111111011110 		: log = 32'b00000000000000001011000001100001;
			12'b111111011111 		: log = 32'b00000000000000001011000001101001;
			12'b111111100000 		: log = 32'b00000000000000001011000001110001;
			12'b111111100001 		: log = 32'b00000000000000001011000001111001;
			12'b111111100010 		: log = 32'b00000000000000001011000010000001;
			12'b111111100011 		: log = 32'b00000000000000001011000010001001;
			12'b111111100100 		: log = 32'b00000000000000001011000010010001;
			12'b111111100101 		: log = 32'b00000000000000001011000010011001;
			12'b111111100110 		: log = 32'b00000000000000001011000010100001;
			12'b111111100111 		: log = 32'b00000000000000001011000010101001;
			12'b111111101000 		: log = 32'b00000000000000001011000010110001;
			12'b111111101001 		: log = 32'b00000000000000001011000010111001;
			12'b111111101010 		: log = 32'b00000000000000001011000011000001;
			12'b111111101011 		: log = 32'b00000000000000001011000011001001;
			12'b111111101100 		: log = 32'b00000000000000001011000011010001;
			12'b111111101101 		: log = 32'b00000000000000001011000011011001;
			12'b111111101110 		: log = 32'b00000000000000001011000011100001;
			12'b111111101111 		: log = 32'b00000000000000001011000011101001;
			12'b111111110000 		: log = 32'b00000000000000001011000011110001;
			12'b111111110001 		: log = 32'b00000000000000001011000011111001;
			12'b111111110010 		: log = 32'b00000000000000001011000100000001;
			12'b111111110011 		: log = 32'b00000000000000001011000100001010;
			12'b111111110100 		: log = 32'b00000000000000001011000100010010;
			12'b111111110101 		: log = 32'b00000000000000001011000100011010;
			12'b111111110110 		: log = 32'b00000000000000001011000100100010;
			12'b111111110111 		: log = 32'b00000000000000001011000100101010;
			12'b111111111000 		: log = 32'b00000000000000001011000100110010;
			12'b111111111001 		: log = 32'b00000000000000001011000100111010;
			12'b111111111010 		: log = 32'b00000000000000001011000101000010;
			12'b111111111011 		: log = 32'b00000000000000001011000101001010;
			12'b111111111100 		: log = 32'b00000000000000001011000101010010;
			12'b111111111101 		: log = 32'b00000000000000001011000101011010;
			12'b111111111110 		: log = 32'b00000000000000001011000101100010;
			12'b111111111111 		: log = 32'b00000000000000001011000101101010;
        endcase
    end
endmodule
