module LUT2(addr, log);
    input [9:0] addr;
    output reg [15:0] log;

    always @(addr) begin
        case (addr)
			10'b0 		: log = 16'b0000000000000000;
			10'b1 		: log = 16'b0001001111111111;
			10'b10 		: log = 16'b0001011111111110;
			10'b11 		: log = 16'b0001100111111110;
			10'b100 		: log = 16'b0001101111111100;
			10'b101 		: log = 16'b0001110011111101;
			10'b110 		: log = 16'b0001110111111100;
			10'b111 		: log = 16'b0001111011111010;
			10'b1000 		: log = 16'b0001111111111000;
			10'b1001 		: log = 16'b0010000001111011;
			10'b1010 		: log = 16'b0010000011111010;
			10'b1011 		: log = 16'b0010000101111000;
			10'b1100 		: log = 16'b0010000111110111;
			10'b1101 		: log = 16'b0010001001110110;
			10'b1110 		: log = 16'b0010001011110100;
			10'b1111 		: log = 16'b0010001101110010;
			10'b10000 		: log = 16'b0010001111110000;
			10'b10001 		: log = 16'b0010010000110111;
			10'b10010 		: log = 16'b0010010001110110;
			10'b10011 		: log = 16'b0010010010110101;
			10'b10100 		: log = 16'b0010010011110100;
			10'b10101 		: log = 16'b0010010100110010;
			10'b10110 		: log = 16'b0010010101110001;
			10'b10111 		: log = 16'b0010010110110000;
			10'b11000 		: log = 16'b0010010111101110;
			10'b11001 		: log = 16'b0010011000101101;
			10'b11010 		: log = 16'b0010011001101011;
			10'b11011 		: log = 16'b0010011010101010;
			10'b11100 		: log = 16'b0010011011101000;
			10'b11101 		: log = 16'b0010011100100110;
			10'b11110 		: log = 16'b0010011101100100;
			10'b11111 		: log = 16'b0010011110100011;
			10'b100000 		: log = 16'b0010011111100001;
			10'b100001 		: log = 16'b0010100000001111;
			10'b100010 		: log = 16'b0010100000101110;
			10'b100011 		: log = 16'b0010100001001101;
			10'b100100 		: log = 16'b0010100001101100;
			10'b100101 		: log = 16'b0010100010001011;
			10'b100110 		: log = 16'b0010100010101010;
			10'b100111 		: log = 16'b0010100011001001;
			10'b101000 		: log = 16'b0010100011101000;
			10'b101001 		: log = 16'b0010100100000110;
			10'b101010 		: log = 16'b0010100100100101;
			10'b101011 		: log = 16'b0010100101000100;
			10'b101100 		: log = 16'b0010100101100011;
			10'b101101 		: log = 16'b0010100110000001;
			10'b101110 		: log = 16'b0010100110100000;
			10'b101111 		: log = 16'b0010100110111111;
			10'b110000 		: log = 16'b0010100111011101;
			10'b110001 		: log = 16'b0010100111111100;
			10'b110010 		: log = 16'b0010101000011010;
			10'b110011 		: log = 16'b0010101000111001;
			10'b110100 		: log = 16'b0010101001010111;
			10'b110101 		: log = 16'b0010101001110110;
			10'b110110 		: log = 16'b0010101010010100;
			10'b110111 		: log = 16'b0010101010110010;
			10'b111000 		: log = 16'b0010101011010001;
			10'b111001 		: log = 16'b0010101011101111;
			10'b111010 		: log = 16'b0010101100001101;
			10'b111011 		: log = 16'b0010101100101100;
			10'b111100 		: log = 16'b0010101101001010;
			10'b111101 		: log = 16'b0010101101101000;
			10'b111110 		: log = 16'b0010101110000110;
			10'b111111 		: log = 16'b0010101110100100;
			10'b1000000 		: log = 16'b0010101111000011;
			10'b1000001 		: log = 16'b0010101111100001;
			10'b1000010 		: log = 16'b0010101111111111;
			10'b1000011 		: log = 16'b0010110000001110;
			10'b1000100 		: log = 16'b0010110000011101;
			10'b1000101 		: log = 16'b0010110000101100;
			10'b1000110 		: log = 16'b0010110000111011;
			10'b1000111 		: log = 16'b0010110001001010;
			10'b1001000 		: log = 16'b0010110001011001;
			10'b1001001 		: log = 16'b0010110001101000;
			10'b1001010 		: log = 16'b0010110001110111;
			10'b1001011 		: log = 16'b0010110010000110;
			10'b1001100 		: log = 16'b0010110010010101;
			10'b1001101 		: log = 16'b0010110010100100;
			10'b1001110 		: log = 16'b0010110010110011;
			10'b1001111 		: log = 16'b0010110011000010;
			10'b1010000 		: log = 16'b0010110011010000;
			10'b1010001 		: log = 16'b0010110011011111;
			10'b1010010 		: log = 16'b0010110011101110;
			10'b1010011 		: log = 16'b0010110011111101;
			10'b1010100 		: log = 16'b0010110100001100;
			10'b1010101 		: log = 16'b0010110100011010;
			10'b1010110 		: log = 16'b0010110100101001;
			10'b1010111 		: log = 16'b0010110100111000;
			10'b1011000 		: log = 16'b0010110101000111;
			10'b1011001 		: log = 16'b0010110101010101;
			10'b1011010 		: log = 16'b0010110101100100;
			10'b1011011 		: log = 16'b0010110101110011;
			10'b1011100 		: log = 16'b0010110110000010;
			10'b1011101 		: log = 16'b0010110110010000;
			10'b1011110 		: log = 16'b0010110110011111;
			10'b1011111 		: log = 16'b0010110110101110;
			10'b1100000 		: log = 16'b0010110110111100;
			10'b1100001 		: log = 16'b0010110111001011;
			10'b1100010 		: log = 16'b0010110111011001;
			10'b1100011 		: log = 16'b0010110111101000;
			10'b1100100 		: log = 16'b0010110111110111;
			10'b1100101 		: log = 16'b0010111000000101;
			10'b1100110 		: log = 16'b0010111000010100;
			10'b1100111 		: log = 16'b0010111000100010;
			10'b1101000 		: log = 16'b0010111000110001;
			10'b1101001 		: log = 16'b0010111000111111;
			10'b1101010 		: log = 16'b0010111001001110;
			10'b1101011 		: log = 16'b0010111001011100;
			10'b1101100 		: log = 16'b0010111001101011;
			10'b1101101 		: log = 16'b0010111001111001;
			10'b1101110 		: log = 16'b0010111010001000;
			10'b1101111 		: log = 16'b0010111010010110;
			10'b1110000 		: log = 16'b0010111010100101;
			10'b1110001 		: log = 16'b0010111010110011;
			10'b1110010 		: log = 16'b0010111011000001;
			10'b1110011 		: log = 16'b0010111011010000;
			10'b1110100 		: log = 16'b0010111011011110;
			10'b1110101 		: log = 16'b0010111011101101;
			10'b1110110 		: log = 16'b0010111011111011;
			10'b1110111 		: log = 16'b0010111100001001;
			10'b1111000 		: log = 16'b0010111100011000;
			10'b1111001 		: log = 16'b0010111100100110;
			10'b1111010 		: log = 16'b0010111100110100;
			10'b1111011 		: log = 16'b0010111101000010;
			10'b1111100 		: log = 16'b0010111101010001;
			10'b1111101 		: log = 16'b0010111101011111;
			10'b1111110 		: log = 16'b0010111101101101;
			10'b1111111 		: log = 16'b0010111101111100;
			10'b10000000 		: log = 16'b0010111110001010;
			10'b10000001 		: log = 16'b0010111110011000;
			10'b10000010 		: log = 16'b0010111110100110;
			10'b10000011 		: log = 16'b0010111110110100;
			10'b10000100 		: log = 16'b0010111111000011;
			10'b10000101 		: log = 16'b0010111111010001;
			10'b10000110 		: log = 16'b0010111111011111;
			10'b10000111 		: log = 16'b0010111111101101;
			10'b10001000 		: log = 16'b0010111111111011;
			10'b10001001 		: log = 16'b0011000000000101;
			10'b10001010 		: log = 16'b0011000000001100;
			10'b10001011 		: log = 16'b0011000000010011;
			10'b10001100 		: log = 16'b0011000000011010;
			10'b10001101 		: log = 16'b0011000000100001;
			10'b10001110 		: log = 16'b0011000000101000;
			10'b10001111 		: log = 16'b0011000000101111;
			10'b10010000 		: log = 16'b0011000000110110;
			10'b10010001 		: log = 16'b0011000000111101;
			10'b10010010 		: log = 16'b0011000001000100;
			10'b10010011 		: log = 16'b0011000001001011;
			10'b10010100 		: log = 16'b0011000001010010;
			10'b10010101 		: log = 16'b0011000001011001;
			10'b10010110 		: log = 16'b0011000001100000;
			10'b10010111 		: log = 16'b0011000001100111;
			10'b10011000 		: log = 16'b0011000001101110;
			10'b10011001 		: log = 16'b0011000001110101;
			10'b10011010 		: log = 16'b0011000001111100;
			10'b10011011 		: log = 16'b0011000010000011;
			10'b10011100 		: log = 16'b0011000010001010;
			10'b10011101 		: log = 16'b0011000010010001;
			10'b10011110 		: log = 16'b0011000010010111;
			10'b10011111 		: log = 16'b0011000010011110;
			10'b10100000 		: log = 16'b0011000010100101;
			10'b10100001 		: log = 16'b0011000010101100;
			10'b10100010 		: log = 16'b0011000010110011;
			10'b10100011 		: log = 16'b0011000010111010;
			10'b10100100 		: log = 16'b0011000011000001;
			10'b10100101 		: log = 16'b0011000011001000;
			10'b10100110 		: log = 16'b0011000011001111;
			10'b10100111 		: log = 16'b0011000011010110;
			10'b10101000 		: log = 16'b0011000011011100;
			10'b10101001 		: log = 16'b0011000011100011;
			10'b10101010 		: log = 16'b0011000011101010;
			10'b10101011 		: log = 16'b0011000011110001;
			10'b10101100 		: log = 16'b0011000011111000;
			10'b10101101 		: log = 16'b0011000011111111;
			10'b10101110 		: log = 16'b0011000100000110;
			10'b10101111 		: log = 16'b0011000100001100;
			10'b10110000 		: log = 16'b0011000100010011;
			10'b10110001 		: log = 16'b0011000100011010;
			10'b10110010 		: log = 16'b0011000100100001;
			10'b10110011 		: log = 16'b0011000100101000;
			10'b10110100 		: log = 16'b0011000100101111;
			10'b10110101 		: log = 16'b0011000100110101;
			10'b10110110 		: log = 16'b0011000100111100;
			10'b10110111 		: log = 16'b0011000101000011;
			10'b10111000 		: log = 16'b0011000101001010;
			10'b10111001 		: log = 16'b0011000101010001;
			10'b10111010 		: log = 16'b0011000101010111;
			10'b10111011 		: log = 16'b0011000101011110;
			10'b10111100 		: log = 16'b0011000101100101;
			10'b10111101 		: log = 16'b0011000101101100;
			10'b10111110 		: log = 16'b0011000101110010;
			10'b10111111 		: log = 16'b0011000101111001;
			10'b11000000 		: log = 16'b0011000110000000;
			10'b11000001 		: log = 16'b0011000110000111;
			10'b11000010 		: log = 16'b0011000110001101;
			10'b11000011 		: log = 16'b0011000110010100;
			10'b11000100 		: log = 16'b0011000110011011;
			10'b11000101 		: log = 16'b0011000110100001;
			10'b11000110 		: log = 16'b0011000110101000;
			10'b11000111 		: log = 16'b0011000110101111;
			10'b11001000 		: log = 16'b0011000110110110;
			10'b11001001 		: log = 16'b0011000110111100;
			10'b11001010 		: log = 16'b0011000111000011;
			10'b11001011 		: log = 16'b0011000111001010;
			10'b11001100 		: log = 16'b0011000111010000;
			10'b11001101 		: log = 16'b0011000111010111;
			10'b11001110 		: log = 16'b0011000111011110;
			10'b11001111 		: log = 16'b0011000111100100;
			10'b11010000 		: log = 16'b0011000111101011;
			10'b11010001 		: log = 16'b0011000111110010;
			10'b11010010 		: log = 16'b0011000111111000;
			10'b11010011 		: log = 16'b0011000111111111;
			10'b11010100 		: log = 16'b0011001000000101;
			10'b11010101 		: log = 16'b0011001000001100;
			10'b11010110 		: log = 16'b0011001000010011;
			10'b11010111 		: log = 16'b0011001000011001;
			10'b11011000 		: log = 16'b0011001000100000;
			10'b11011001 		: log = 16'b0011001000100111;
			10'b11011010 		: log = 16'b0011001000101101;
			10'b11011011 		: log = 16'b0011001000110100;
			10'b11011100 		: log = 16'b0011001000111010;
			10'b11011101 		: log = 16'b0011001001000001;
			10'b11011110 		: log = 16'b0011001001000111;
			10'b11011111 		: log = 16'b0011001001001110;
			10'b11100000 		: log = 16'b0011001001010101;
			10'b11100001 		: log = 16'b0011001001011011;
			10'b11100010 		: log = 16'b0011001001100010;
			10'b11100011 		: log = 16'b0011001001101000;
			10'b11100100 		: log = 16'b0011001001101111;
			10'b11100101 		: log = 16'b0011001001110101;
			10'b11100110 		: log = 16'b0011001001111100;
			10'b11100111 		: log = 16'b0011001010000010;
			10'b11101000 		: log = 16'b0011001010001001;
			10'b11101001 		: log = 16'b0011001010001111;
			10'b11101010 		: log = 16'b0011001010010110;
			10'b11101011 		: log = 16'b0011001010011100;
			10'b11101100 		: log = 16'b0011001010100011;
			10'b11101101 		: log = 16'b0011001010101001;
			10'b11101110 		: log = 16'b0011001010110000;
			10'b11101111 		: log = 16'b0011001010110110;
			10'b11110000 		: log = 16'b0011001010111101;
			10'b11110001 		: log = 16'b0011001011000011;
			10'b11110010 		: log = 16'b0011001011001010;
			10'b11110011 		: log = 16'b0011001011010000;
			10'b11110100 		: log = 16'b0011001011010111;
			10'b11110101 		: log = 16'b0011001011011101;
			10'b11110110 		: log = 16'b0011001011100100;
			10'b11110111 		: log = 16'b0011001011101010;
			10'b11111000 		: log = 16'b0011001011110001;
			10'b11111001 		: log = 16'b0011001011110111;
			10'b11111010 		: log = 16'b0011001011111110;
			10'b11111011 		: log = 16'b0011001100000100;
			10'b11111100 		: log = 16'b0011001100001010;
			10'b11111101 		: log = 16'b0011001100010001;
			10'b11111110 		: log = 16'b0011001100010111;
			10'b11111111 		: log = 16'b0011001100011110;
			10'b100000000 		: log = 16'b0011001100100100;
			10'b100000001 		: log = 16'b0011001100101010;
			10'b100000010 		: log = 16'b0011001100110001;
			10'b100000011 		: log = 16'b0011001100110111;
			10'b100000100 		: log = 16'b0011001100111110;
			10'b100000101 		: log = 16'b0011001101000100;
			10'b100000110 		: log = 16'b0011001101001010;
			10'b100000111 		: log = 16'b0011001101010001;
			10'b100001000 		: log = 16'b0011001101010111;
			10'b100001001 		: log = 16'b0011001101011101;
			10'b100001010 		: log = 16'b0011001101100100;
			10'b100001011 		: log = 16'b0011001101101010;
			10'b100001100 		: log = 16'b0011001101110000;
			10'b100001101 		: log = 16'b0011001101110111;
			10'b100001110 		: log = 16'b0011001101111101;
			10'b100001111 		: log = 16'b0011001110000011;
			10'b100010000 		: log = 16'b0011001110001010;
			10'b100010001 		: log = 16'b0011001110010000;
			10'b100010010 		: log = 16'b0011001110010110;
			10'b100010011 		: log = 16'b0011001110011101;
			10'b100010100 		: log = 16'b0011001110100011;
			10'b100010101 		: log = 16'b0011001110101001;
			10'b100010110 		: log = 16'b0011001110110000;
			10'b100010111 		: log = 16'b0011001110110110;
			10'b100011000 		: log = 16'b0011001110111100;
			10'b100011001 		: log = 16'b0011001111000010;
			10'b100011010 		: log = 16'b0011001111001001;
			10'b100011011 		: log = 16'b0011001111001111;
			10'b100011100 		: log = 16'b0011001111010101;
			10'b100011101 		: log = 16'b0011001111011100;
			10'b100011110 		: log = 16'b0011001111100010;
			10'b100011111 		: log = 16'b0011001111101000;
			10'b100100000 		: log = 16'b0011001111101110;
			10'b100100001 		: log = 16'b0011001111110101;
			10'b100100010 		: log = 16'b0011001111111011;
			10'b100100011 		: log = 16'b0011010000000000;
			10'b100100100 		: log = 16'b0011010000000100;
			10'b100100101 		: log = 16'b0011010000000111;
			10'b100100110 		: log = 16'b0011010000001010;
			10'b100100111 		: log = 16'b0011010000001101;
			10'b100101000 		: log = 16'b0011010000010000;
			10'b100101001 		: log = 16'b0011010000010011;
			10'b100101010 		: log = 16'b0011010000010110;
			10'b100101011 		: log = 16'b0011010000011001;
			10'b100101100 		: log = 16'b0011010000011100;
			10'b100101101 		: log = 16'b0011010000100000;
			10'b100101110 		: log = 16'b0011010000100011;
			10'b100101111 		: log = 16'b0011010000100110;
			10'b100110000 		: log = 16'b0011010000101001;
			10'b100110001 		: log = 16'b0011010000101100;
			10'b100110010 		: log = 16'b0011010000101111;
			10'b100110011 		: log = 16'b0011010000110010;
			10'b100110100 		: log = 16'b0011010000110101;
			10'b100110101 		: log = 16'b0011010000111000;
			10'b100110110 		: log = 16'b0011010000111011;
			10'b100110111 		: log = 16'b0011010000111110;
			10'b100111000 		: log = 16'b0011010001000001;
			10'b100111001 		: log = 16'b0011010001000100;
			10'b100111010 		: log = 16'b0011010001001000;
			10'b100111011 		: log = 16'b0011010001001011;
			10'b100111100 		: log = 16'b0011010001001110;
			10'b100111101 		: log = 16'b0011010001010001;
			10'b100111110 		: log = 16'b0011010001010100;
			10'b100111111 		: log = 16'b0011010001010111;
			10'b101000000 		: log = 16'b0011010001011010;
			10'b101000001 		: log = 16'b0011010001011101;
			10'b101000010 		: log = 16'b0011010001100000;
			10'b101000011 		: log = 16'b0011010001100011;
			10'b101000100 		: log = 16'b0011010001100110;
			10'b101000101 		: log = 16'b0011010001101001;
			10'b101000110 		: log = 16'b0011010001101100;
			10'b101000111 		: log = 16'b0011010001101111;
			10'b101001000 		: log = 16'b0011010001110010;
			10'b101001001 		: log = 16'b0011010001110101;
			10'b101001010 		: log = 16'b0011010001111000;
			10'b101001011 		: log = 16'b0011010001111011;
			10'b101001100 		: log = 16'b0011010001111110;
			10'b101001101 		: log = 16'b0011010010000001;
			10'b101001110 		: log = 16'b0011010010000100;
			10'b101001111 		: log = 16'b0011010010000111;
			10'b101010000 		: log = 16'b0011010010001010;
			10'b101010001 		: log = 16'b0011010010001101;
			10'b101010010 		: log = 16'b0011010010010000;
			10'b101010011 		: log = 16'b0011010010010011;
			10'b101010100 		: log = 16'b0011010010010110;
			10'b101010101 		: log = 16'b0011010010011001;
			10'b101010110 		: log = 16'b0011010010011100;
			10'b101010111 		: log = 16'b0011010010011111;
			10'b101011000 		: log = 16'b0011010010100010;
			10'b101011001 		: log = 16'b0011010010100101;
			10'b101011010 		: log = 16'b0011010010101000;
			10'b101011011 		: log = 16'b0011010010101011;
			10'b101011100 		: log = 16'b0011010010101110;
			10'b101011101 		: log = 16'b0011010010110001;
			10'b101011110 		: log = 16'b0011010010110100;
			10'b101011111 		: log = 16'b0011010010110111;
			10'b101100000 		: log = 16'b0011010010111010;
			10'b101100001 		: log = 16'b0011010010111101;
			10'b101100010 		: log = 16'b0011010011000000;
			10'b101100011 		: log = 16'b0011010011000011;
			10'b101100100 		: log = 16'b0011010011000110;
			10'b101100101 		: log = 16'b0011010011001001;
			10'b101100110 		: log = 16'b0011010011001100;
			10'b101100111 		: log = 16'b0011010011001111;
			10'b101101000 		: log = 16'b0011010011010010;
			10'b101101001 		: log = 16'b0011010011010101;
			10'b101101010 		: log = 16'b0011010011011000;
			10'b101101011 		: log = 16'b0011010011011011;
			10'b101101100 		: log = 16'b0011010011011110;
			10'b101101101 		: log = 16'b0011010011100001;
			10'b101101110 		: log = 16'b0011010011100100;
			10'b101101111 		: log = 16'b0011010011100111;
			10'b101110000 		: log = 16'b0011010011101010;
			10'b101110001 		: log = 16'b0011010011101101;
			10'b101110010 		: log = 16'b0011010011101111;
			10'b101110011 		: log = 16'b0011010011110010;
			10'b101110100 		: log = 16'b0011010011110101;
			10'b101110101 		: log = 16'b0011010011111000;
			10'b101110110 		: log = 16'b0011010011111011;
			10'b101110111 		: log = 16'b0011010011111110;
			10'b101111000 		: log = 16'b0011010100000001;
			10'b101111001 		: log = 16'b0011010100000100;
			10'b101111010 		: log = 16'b0011010100000111;
			10'b101111011 		: log = 16'b0011010100001010;
			10'b101111100 		: log = 16'b0011010100001101;
			10'b101111101 		: log = 16'b0011010100010000;
			10'b101111110 		: log = 16'b0011010100010011;
			10'b101111111 		: log = 16'b0011010100010101;
			10'b110000000 		: log = 16'b0011010100011000;
			10'b110000001 		: log = 16'b0011010100011011;
			10'b110000010 		: log = 16'b0011010100011110;
			10'b110000011 		: log = 16'b0011010100100001;
			10'b110000100 		: log = 16'b0011010100100100;
			10'b110000101 		: log = 16'b0011010100100111;
			10'b110000110 		: log = 16'b0011010100101010;
			10'b110000111 		: log = 16'b0011010100101101;
			10'b110001000 		: log = 16'b0011010100110000;
			10'b110001001 		: log = 16'b0011010100110010;
			10'b110001010 		: log = 16'b0011010100110101;
			10'b110001011 		: log = 16'b0011010100111000;
			10'b110001100 		: log = 16'b0011010100111011;
			10'b110001101 		: log = 16'b0011010100111110;
			10'b110001110 		: log = 16'b0011010101000001;
			10'b110001111 		: log = 16'b0011010101000100;
			10'b110010000 		: log = 16'b0011010101000111;
			10'b110010001 		: log = 16'b0011010101001010;
			10'b110010010 		: log = 16'b0011010101001100;
			10'b110010011 		: log = 16'b0011010101001111;
			10'b110010100 		: log = 16'b0011010101010010;
			10'b110010101 		: log = 16'b0011010101010101;
			10'b110010110 		: log = 16'b0011010101011000;
			10'b110010111 		: log = 16'b0011010101011011;
			10'b110011000 		: log = 16'b0011010101011110;
			10'b110011001 		: log = 16'b0011010101100000;
			10'b110011010 		: log = 16'b0011010101100011;
			10'b110011011 		: log = 16'b0011010101100110;
			10'b110011100 		: log = 16'b0011010101101001;
			10'b110011101 		: log = 16'b0011010101101100;
			10'b110011110 		: log = 16'b0011010101101111;
			10'b110011111 		: log = 16'b0011010101110010;
			10'b110100000 		: log = 16'b0011010101110100;
			10'b110100001 		: log = 16'b0011010101110111;
			10'b110100010 		: log = 16'b0011010101111010;
			10'b110100011 		: log = 16'b0011010101111101;
			10'b110100100 		: log = 16'b0011010110000000;
			10'b110100101 		: log = 16'b0011010110000011;
			10'b110100110 		: log = 16'b0011010110000101;
			10'b110100111 		: log = 16'b0011010110001000;
			10'b110101000 		: log = 16'b0011010110001011;
			10'b110101001 		: log = 16'b0011010110001110;
			10'b110101010 		: log = 16'b0011010110010001;
			10'b110101011 		: log = 16'b0011010110010100;
			10'b110101100 		: log = 16'b0011010110010110;
			10'b110101101 		: log = 16'b0011010110011001;
			10'b110101110 		: log = 16'b0011010110011100;
			10'b110101111 		: log = 16'b0011010110011111;
			10'b110110000 		: log = 16'b0011010110100010;
			10'b110110001 		: log = 16'b0011010110100101;
			10'b110110010 		: log = 16'b0011010110100111;
			10'b110110011 		: log = 16'b0011010110101010;
			10'b110110100 		: log = 16'b0011010110101101;
			10'b110110101 		: log = 16'b0011010110110000;
			10'b110110110 		: log = 16'b0011010110110011;
			10'b110110111 		: log = 16'b0011010110110101;
			10'b110111000 		: log = 16'b0011010110111000;
			10'b110111001 		: log = 16'b0011010110111011;
			10'b110111010 		: log = 16'b0011010110111110;
			10'b110111011 		: log = 16'b0011010111000001;
			10'b110111100 		: log = 16'b0011010111000011;
			10'b110111101 		: log = 16'b0011010111000110;
			10'b110111110 		: log = 16'b0011010111001001;
			10'b110111111 		: log = 16'b0011010111001100;
			10'b111000000 		: log = 16'b0011010111001110;
			10'b111000001 		: log = 16'b0011010111010001;
			10'b111000010 		: log = 16'b0011010111010100;
			10'b111000011 		: log = 16'b0011010111010111;
			10'b111000100 		: log = 16'b0011010111011010;
			10'b111000101 		: log = 16'b0011010111011100;
			10'b111000110 		: log = 16'b0011010111011111;
			10'b111000111 		: log = 16'b0011010111100010;
			10'b111001000 		: log = 16'b0011010111100101;
			10'b111001001 		: log = 16'b0011010111100111;
			10'b111001010 		: log = 16'b0011010111101010;
			10'b111001011 		: log = 16'b0011010111101101;
			10'b111001100 		: log = 16'b0011010111110000;
			10'b111001101 		: log = 16'b0011010111110010;
			10'b111001110 		: log = 16'b0011010111110101;
			10'b111001111 		: log = 16'b0011010111111000;
			10'b111010000 		: log = 16'b0011010111111011;
			10'b111010001 		: log = 16'b0011010111111101;
			10'b111010010 		: log = 16'b0011011000000000;
			10'b111010011 		: log = 16'b0011011000000011;
			10'b111010100 		: log = 16'b0011011000000110;
			10'b111010101 		: log = 16'b0011011000001000;
			10'b111010110 		: log = 16'b0011011000001011;
			10'b111010111 		: log = 16'b0011011000001110;
			10'b111011000 		: log = 16'b0011011000010001;
			10'b111011001 		: log = 16'b0011011000010011;
			10'b111011010 		: log = 16'b0011011000010110;
			10'b111011011 		: log = 16'b0011011000011001;
			10'b111011100 		: log = 16'b0011011000011100;
			10'b111011101 		: log = 16'b0011011000011110;
			10'b111011110 		: log = 16'b0011011000100001;
			10'b111011111 		: log = 16'b0011011000100100;
			10'b111100000 		: log = 16'b0011011000100111;
			10'b111100001 		: log = 16'b0011011000101001;
			10'b111100010 		: log = 16'b0011011000101100;
			10'b111100011 		: log = 16'b0011011000101111;
			10'b111100100 		: log = 16'b0011011000110001;
			10'b111100101 		: log = 16'b0011011000110100;
			10'b111100110 		: log = 16'b0011011000110111;
			10'b111100111 		: log = 16'b0011011000111010;
			10'b111101000 		: log = 16'b0011011000111100;
			10'b111101001 		: log = 16'b0011011000111111;
			10'b111101010 		: log = 16'b0011011001000010;
			10'b111101011 		: log = 16'b0011011001000100;
			10'b111101100 		: log = 16'b0011011001000111;
			10'b111101101 		: log = 16'b0011011001001010;
			10'b111101110 		: log = 16'b0011011001001101;
			10'b111101111 		: log = 16'b0011011001001111;
			10'b111110000 		: log = 16'b0011011001010010;
			10'b111110001 		: log = 16'b0011011001010101;
			10'b111110010 		: log = 16'b0011011001010111;
			10'b111110011 		: log = 16'b0011011001011010;
			10'b111110100 		: log = 16'b0011011001011101;
			10'b111110101 		: log = 16'b0011011001011111;
			10'b111110110 		: log = 16'b0011011001100010;
			10'b111110111 		: log = 16'b0011011001100101;
			10'b111111000 		: log = 16'b0011011001100111;
			10'b111111001 		: log = 16'b0011011001101010;
			10'b111111010 		: log = 16'b0011011001101101;
			10'b111111011 		: log = 16'b0011011001101111;
			10'b111111100 		: log = 16'b0011011001110010;
			10'b111111101 		: log = 16'b0011011001110101;
			10'b111111110 		: log = 16'b0011011001110111;
			10'b111111111 		: log = 16'b0011011001111010;
			10'b1000000000 		: log = 16'b0011011001111101;
			10'b1000000001 		: log = 16'b0011011001111111;
			10'b1000000010 		: log = 16'b0011011010000010;
			10'b1000000011 		: log = 16'b0011011010000101;
			10'b1000000100 		: log = 16'b0011011010000111;
			10'b1000000101 		: log = 16'b0011011010001010;
			10'b1000000110 		: log = 16'b0011011010001101;
			10'b1000000111 		: log = 16'b0011011010001111;
			10'b1000001000 		: log = 16'b0011011010010010;
			10'b1000001001 		: log = 16'b0011011010010101;
			10'b1000001010 		: log = 16'b0011011010010111;
			10'b1000001011 		: log = 16'b0011011010011010;
			10'b1000001100 		: log = 16'b0011011010011101;
			10'b1000001101 		: log = 16'b0011011010011111;
			10'b1000001110 		: log = 16'b0011011010100010;
			10'b1000001111 		: log = 16'b0011011010100101;
			10'b1000010000 		: log = 16'b0011011010100111;
			10'b1000010001 		: log = 16'b0011011010101010;
			10'b1000010010 		: log = 16'b0011011010101101;
			10'b1000010011 		: log = 16'b0011011010101111;
			10'b1000010100 		: log = 16'b0011011010110010;
			10'b1000010101 		: log = 16'b0011011010110100;
			10'b1000010110 		: log = 16'b0011011010110111;
			10'b1000010111 		: log = 16'b0011011010111010;
			10'b1000011000 		: log = 16'b0011011010111100;
			10'b1000011001 		: log = 16'b0011011010111111;
			10'b1000011010 		: log = 16'b0011011011000010;
			10'b1000011011 		: log = 16'b0011011011000100;
			10'b1000011100 		: log = 16'b0011011011000111;
			10'b1000011101 		: log = 16'b0011011011001001;
			10'b1000011110 		: log = 16'b0011011011001100;
			10'b1000011111 		: log = 16'b0011011011001111;
			10'b1000100000 		: log = 16'b0011011011010001;
			10'b1000100001 		: log = 16'b0011011011010100;
			10'b1000100010 		: log = 16'b0011011011010110;
			10'b1000100011 		: log = 16'b0011011011011001;
			10'b1000100100 		: log = 16'b0011011011011100;
			10'b1000100101 		: log = 16'b0011011011011110;
			10'b1000100110 		: log = 16'b0011011011100001;
			10'b1000100111 		: log = 16'b0011011011100011;
			10'b1000101000 		: log = 16'b0011011011100110;
			10'b1000101001 		: log = 16'b0011011011101001;
			10'b1000101010 		: log = 16'b0011011011101011;
			10'b1000101011 		: log = 16'b0011011011101110;
			10'b1000101100 		: log = 16'b0011011011110000;
			10'b1000101101 		: log = 16'b0011011011110011;
			10'b1000101110 		: log = 16'b0011011011110110;
			10'b1000101111 		: log = 16'b0011011011111000;
			10'b1000110000 		: log = 16'b0011011011111011;
			10'b1000110001 		: log = 16'b0011011011111101;
			10'b1000110010 		: log = 16'b0011011100000000;
			10'b1000110011 		: log = 16'b0011011100000011;
			10'b1000110100 		: log = 16'b0011011100000101;
			10'b1000110101 		: log = 16'b0011011100001000;
			10'b1000110110 		: log = 16'b0011011100001010;
			10'b1000110111 		: log = 16'b0011011100001101;
			10'b1000111000 		: log = 16'b0011011100001111;
			10'b1000111001 		: log = 16'b0011011100010010;
			10'b1000111010 		: log = 16'b0011011100010101;
			10'b1000111011 		: log = 16'b0011011100010111;
			10'b1000111100 		: log = 16'b0011011100011010;
			10'b1000111101 		: log = 16'b0011011100011100;
			10'b1000111110 		: log = 16'b0011011100011111;
			10'b1000111111 		: log = 16'b0011011100100001;
			10'b1001000000 		: log = 16'b0011011100100100;
			10'b1001000001 		: log = 16'b0011011100100111;
			10'b1001000010 		: log = 16'b0011011100101001;
			10'b1001000011 		: log = 16'b0011011100101100;
			10'b1001000100 		: log = 16'b0011011100101110;
			10'b1001000101 		: log = 16'b0011011100110001;
			10'b1001000110 		: log = 16'b0011011100110011;
			10'b1001000111 		: log = 16'b0011011100110110;
			10'b1001001000 		: log = 16'b0011011100111000;
			10'b1001001001 		: log = 16'b0011011100111011;
			10'b1001001010 		: log = 16'b0011011100111110;
			10'b1001001011 		: log = 16'b0011011101000000;
			10'b1001001100 		: log = 16'b0011011101000011;
			10'b1001001101 		: log = 16'b0011011101000101;
			10'b1001001110 		: log = 16'b0011011101001000;
			10'b1001001111 		: log = 16'b0011011101001010;
			10'b1001010000 		: log = 16'b0011011101001101;
			10'b1001010001 		: log = 16'b0011011101001111;
			10'b1001010010 		: log = 16'b0011011101010010;
			10'b1001010011 		: log = 16'b0011011101010100;
			10'b1001010100 		: log = 16'b0011011101010111;
			10'b1001010101 		: log = 16'b0011011101011001;
			10'b1001010110 		: log = 16'b0011011101011100;
			10'b1001010111 		: log = 16'b0011011101011110;
			10'b1001011000 		: log = 16'b0011011101100001;
			10'b1001011001 		: log = 16'b0011011101100011;
			10'b1001011010 		: log = 16'b0011011101100110;
			10'b1001011011 		: log = 16'b0011011101101001;
			10'b1001011100 		: log = 16'b0011011101101011;
			10'b1001011101 		: log = 16'b0011011101101110;
			10'b1001011110 		: log = 16'b0011011101110000;
			10'b1001011111 		: log = 16'b0011011101110011;
			10'b1001100000 		: log = 16'b0011011101110101;
			10'b1001100001 		: log = 16'b0011011101111000;
			10'b1001100010 		: log = 16'b0011011101111010;
			10'b1001100011 		: log = 16'b0011011101111101;
			10'b1001100100 		: log = 16'b0011011101111111;
			10'b1001100101 		: log = 16'b0011011110000010;
			10'b1001100110 		: log = 16'b0011011110000100;
			10'b1001100111 		: log = 16'b0011011110000111;
			10'b1001101000 		: log = 16'b0011011110001001;
			10'b1001101001 		: log = 16'b0011011110001100;
			10'b1001101010 		: log = 16'b0011011110001110;
			10'b1001101011 		: log = 16'b0011011110010001;
			10'b1001101100 		: log = 16'b0011011110010011;
			10'b1001101101 		: log = 16'b0011011110010110;
			10'b1001101110 		: log = 16'b0011011110011000;
			10'b1001101111 		: log = 16'b0011011110011011;
			10'b1001110000 		: log = 16'b0011011110011101;
			10'b1001110001 		: log = 16'b0011011110100000;
			10'b1001110010 		: log = 16'b0011011110100010;
			10'b1001110011 		: log = 16'b0011011110100101;
			10'b1001110100 		: log = 16'b0011011110100111;
			10'b1001110101 		: log = 16'b0011011110101001;
			10'b1001110110 		: log = 16'b0011011110101100;
			10'b1001110111 		: log = 16'b0011011110101110;
			10'b1001111000 		: log = 16'b0011011110110001;
			10'b1001111001 		: log = 16'b0011011110110011;
			10'b1001111010 		: log = 16'b0011011110110110;
			10'b1001111011 		: log = 16'b0011011110111000;
			10'b1001111100 		: log = 16'b0011011110111011;
			10'b1001111101 		: log = 16'b0011011110111101;
			10'b1001111110 		: log = 16'b0011011111000000;
			10'b1001111111 		: log = 16'b0011011111000010;
			10'b1010000000 		: log = 16'b0011011111000101;
			10'b1010000001 		: log = 16'b0011011111000111;
			10'b1010000010 		: log = 16'b0011011111001010;
			10'b1010000011 		: log = 16'b0011011111001100;
			10'b1010000100 		: log = 16'b0011011111001110;
			10'b1010000101 		: log = 16'b0011011111010001;
			10'b1010000110 		: log = 16'b0011011111010011;
			10'b1010000111 		: log = 16'b0011011111010110;
			10'b1010001000 		: log = 16'b0011011111011000;
			10'b1010001001 		: log = 16'b0011011111011011;
			10'b1010001010 		: log = 16'b0011011111011101;
			10'b1010001011 		: log = 16'b0011011111100000;
			10'b1010001100 		: log = 16'b0011011111100010;
			10'b1010001101 		: log = 16'b0011011111100101;
			10'b1010001110 		: log = 16'b0011011111100111;
			10'b1010001111 		: log = 16'b0011011111101001;
			10'b1010010000 		: log = 16'b0011011111101100;
			10'b1010010001 		: log = 16'b0011011111101110;
			10'b1010010010 		: log = 16'b0011011111110001;
			10'b1010010011 		: log = 16'b0011011111110011;
			10'b1010010100 		: log = 16'b0011011111110110;
			10'b1010010101 		: log = 16'b0011011111111000;
			10'b1010010110 		: log = 16'b0011011111111010;
			10'b1010010111 		: log = 16'b0011011111111101;
			10'b1010011000 		: log = 16'b0011011111111111;
			10'b1010011001 		: log = 16'b0011100000000001;
			10'b1010011010 		: log = 16'b0011100000000010;
			10'b1010011011 		: log = 16'b0011100000000011;
			10'b1010011100 		: log = 16'b0011100000000100;
			10'b1010011101 		: log = 16'b0011100000000110;
			10'b1010011110 		: log = 16'b0011100000000111;
			10'b1010011111 		: log = 16'b0011100000001000;
			10'b1010100000 		: log = 16'b0011100000001001;
			10'b1010100001 		: log = 16'b0011100000001011;
			10'b1010100010 		: log = 16'b0011100000001100;
			10'b1010100011 		: log = 16'b0011100000001101;
			10'b1010100100 		: log = 16'b0011100000001110;
			10'b1010100101 		: log = 16'b0011100000001111;
			10'b1010100110 		: log = 16'b0011100000010001;
			10'b1010100111 		: log = 16'b0011100000010010;
			10'b1010101000 		: log = 16'b0011100000010011;
			10'b1010101001 		: log = 16'b0011100000010100;
			10'b1010101010 		: log = 16'b0011100000010101;
			10'b1010101011 		: log = 16'b0011100000010111;
			10'b1010101100 		: log = 16'b0011100000011000;
			10'b1010101101 		: log = 16'b0011100000011001;
			10'b1010101110 		: log = 16'b0011100000011010;
			10'b1010101111 		: log = 16'b0011100000011011;
			10'b1010110000 		: log = 16'b0011100000011101;
			10'b1010110001 		: log = 16'b0011100000011110;
			10'b1010110010 		: log = 16'b0011100000011111;
			10'b1010110011 		: log = 16'b0011100000100000;
			10'b1010110100 		: log = 16'b0011100000100001;
			10'b1010110101 		: log = 16'b0011100000100011;
			10'b1010110110 		: log = 16'b0011100000100100;
			10'b1010110111 		: log = 16'b0011100000100101;
			10'b1010111000 		: log = 16'b0011100000100110;
			10'b1010111001 		: log = 16'b0011100000100111;
			10'b1010111010 		: log = 16'b0011100000101000;
			10'b1010111011 		: log = 16'b0011100000101010;
			10'b1010111100 		: log = 16'b0011100000101011;
			10'b1010111101 		: log = 16'b0011100000101100;
			10'b1010111110 		: log = 16'b0011100000101101;
			10'b1010111111 		: log = 16'b0011100000101110;
			10'b1011000000 		: log = 16'b0011100000110000;
			10'b1011000001 		: log = 16'b0011100000110001;
			10'b1011000010 		: log = 16'b0011100000110010;
			10'b1011000011 		: log = 16'b0011100000110011;
			10'b1011000100 		: log = 16'b0011100000110100;
			10'b1011000101 		: log = 16'b0011100000110110;
			10'b1011000110 		: log = 16'b0011100000110111;
			10'b1011000111 		: log = 16'b0011100000111000;
			10'b1011001000 		: log = 16'b0011100000111001;
			10'b1011001001 		: log = 16'b0011100000111010;
			10'b1011001010 		: log = 16'b0011100000111011;
			10'b1011001011 		: log = 16'b0011100000111101;
			10'b1011001100 		: log = 16'b0011100000111110;
			10'b1011001101 		: log = 16'b0011100000111111;
			10'b1011001110 		: log = 16'b0011100001000000;
			10'b1011001111 		: log = 16'b0011100001000001;
			10'b1011010000 		: log = 16'b0011100001000010;
			10'b1011010001 		: log = 16'b0011100001000100;
			10'b1011010010 		: log = 16'b0011100001000101;
			10'b1011010011 		: log = 16'b0011100001000110;
			10'b1011010100 		: log = 16'b0011100001000111;
			10'b1011010101 		: log = 16'b0011100001001000;
			10'b1011010110 		: log = 16'b0011100001001010;
			10'b1011010111 		: log = 16'b0011100001001011;
			10'b1011011000 		: log = 16'b0011100001001100;
			10'b1011011001 		: log = 16'b0011100001001101;
			10'b1011011010 		: log = 16'b0011100001001110;
			10'b1011011011 		: log = 16'b0011100001001111;
			10'b1011011100 		: log = 16'b0011100001010001;
			10'b1011011101 		: log = 16'b0011100001010010;
			10'b1011011110 		: log = 16'b0011100001010011;
			10'b1011011111 		: log = 16'b0011100001010100;
			10'b1011100000 		: log = 16'b0011100001010101;
			10'b1011100001 		: log = 16'b0011100001010110;
			10'b1011100010 		: log = 16'b0011100001011000;
			10'b1011100011 		: log = 16'b0011100001011001;
			10'b1011100100 		: log = 16'b0011100001011010;
			10'b1011100101 		: log = 16'b0011100001011011;
			10'b1011100110 		: log = 16'b0011100001011100;
			10'b1011100111 		: log = 16'b0011100001011101;
			10'b1011101000 		: log = 16'b0011100001011110;
			10'b1011101001 		: log = 16'b0011100001100000;
			10'b1011101010 		: log = 16'b0011100001100001;
			10'b1011101011 		: log = 16'b0011100001100010;
			10'b1011101100 		: log = 16'b0011100001100011;
			10'b1011101101 		: log = 16'b0011100001100100;
			10'b1011101110 		: log = 16'b0011100001100101;
			10'b1011101111 		: log = 16'b0011100001100111;
			10'b1011110000 		: log = 16'b0011100001101000;
			10'b1011110001 		: log = 16'b0011100001101001;
			10'b1011110010 		: log = 16'b0011100001101010;
			10'b1011110011 		: log = 16'b0011100001101011;
			10'b1011110100 		: log = 16'b0011100001101100;
			10'b1011110101 		: log = 16'b0011100001101101;
			10'b1011110110 		: log = 16'b0011100001101111;
			10'b1011110111 		: log = 16'b0011100001110000;
			10'b1011111000 		: log = 16'b0011100001110001;
			10'b1011111001 		: log = 16'b0011100001110010;
			10'b1011111010 		: log = 16'b0011100001110011;
			10'b1011111011 		: log = 16'b0011100001110100;
			10'b1011111100 		: log = 16'b0011100001110110;
			10'b1011111101 		: log = 16'b0011100001110111;
			10'b1011111110 		: log = 16'b0011100001111000;
			10'b1011111111 		: log = 16'b0011100001111001;
			10'b1100000000 		: log = 16'b0011100001111010;
			10'b1100000001 		: log = 16'b0011100001111011;
			10'b1100000010 		: log = 16'b0011100001111100;
			10'b1100000011 		: log = 16'b0011100001111110;
			10'b1100000100 		: log = 16'b0011100001111111;
			10'b1100000101 		: log = 16'b0011100010000000;
			10'b1100000110 		: log = 16'b0011100010000001;
			10'b1100000111 		: log = 16'b0011100010000010;
			10'b1100001000 		: log = 16'b0011100010000011;
			10'b1100001001 		: log = 16'b0011100010000100;
			10'b1100001010 		: log = 16'b0011100010000101;
			10'b1100001011 		: log = 16'b0011100010000111;
			10'b1100001100 		: log = 16'b0011100010001000;
			10'b1100001101 		: log = 16'b0011100010001001;
			10'b1100001110 		: log = 16'b0011100010001010;
			10'b1100001111 		: log = 16'b0011100010001011;
			10'b1100010000 		: log = 16'b0011100010001100;
			10'b1100010001 		: log = 16'b0011100010001101;
			10'b1100010010 		: log = 16'b0011100010001111;
			10'b1100010011 		: log = 16'b0011100010010000;
			10'b1100010100 		: log = 16'b0011100010010001;
			10'b1100010101 		: log = 16'b0011100010010010;
			10'b1100010110 		: log = 16'b0011100010010011;
			10'b1100010111 		: log = 16'b0011100010010100;
			10'b1100011000 		: log = 16'b0011100010010101;
			10'b1100011001 		: log = 16'b0011100010010110;
			10'b1100011010 		: log = 16'b0011100010011000;
			10'b1100011011 		: log = 16'b0011100010011001;
			10'b1100011100 		: log = 16'b0011100010011010;
			10'b1100011101 		: log = 16'b0011100010011011;
			10'b1100011110 		: log = 16'b0011100010011100;
			10'b1100011111 		: log = 16'b0011100010011101;
			10'b1100100000 		: log = 16'b0011100010011110;
			10'b1100100001 		: log = 16'b0011100010011111;
			10'b1100100010 		: log = 16'b0011100010100001;
			10'b1100100011 		: log = 16'b0011100010100010;
			10'b1100100100 		: log = 16'b0011100010100011;
			10'b1100100101 		: log = 16'b0011100010100100;
			10'b1100100110 		: log = 16'b0011100010100101;
			10'b1100100111 		: log = 16'b0011100010100110;
			10'b1100101000 		: log = 16'b0011100010100111;
			10'b1100101001 		: log = 16'b0011100010101000;
			10'b1100101010 		: log = 16'b0011100010101010;
			10'b1100101011 		: log = 16'b0011100010101011;
			10'b1100101100 		: log = 16'b0011100010101100;
			10'b1100101101 		: log = 16'b0011100010101101;
			10'b1100101110 		: log = 16'b0011100010101110;
			10'b1100101111 		: log = 16'b0011100010101111;
			10'b1100110000 		: log = 16'b0011100010110000;
			10'b1100110001 		: log = 16'b0011100010110001;
			10'b1100110010 		: log = 16'b0011100010110010;
			10'b1100110011 		: log = 16'b0011100010110100;
			10'b1100110100 		: log = 16'b0011100010110101;
			10'b1100110101 		: log = 16'b0011100010110110;
			10'b1100110110 		: log = 16'b0011100010110111;
			10'b1100110111 		: log = 16'b0011100010111000;
			10'b1100111000 		: log = 16'b0011100010111001;
			10'b1100111001 		: log = 16'b0011100010111010;
			10'b1100111010 		: log = 16'b0011100010111011;
			10'b1100111011 		: log = 16'b0011100010111100;
			10'b1100111100 		: log = 16'b0011100010111110;
			10'b1100111101 		: log = 16'b0011100010111111;
			10'b1100111110 		: log = 16'b0011100011000000;
			10'b1100111111 		: log = 16'b0011100011000001;
			10'b1101000000 		: log = 16'b0011100011000010;
			10'b1101000001 		: log = 16'b0011100011000011;
			10'b1101000010 		: log = 16'b0011100011000100;
			10'b1101000011 		: log = 16'b0011100011000101;
			10'b1101000100 		: log = 16'b0011100011000110;
			10'b1101000101 		: log = 16'b0011100011000111;
			10'b1101000110 		: log = 16'b0011100011001001;
			10'b1101000111 		: log = 16'b0011100011001010;
			10'b1101001000 		: log = 16'b0011100011001011;
			10'b1101001001 		: log = 16'b0011100011001100;
			10'b1101001010 		: log = 16'b0011100011001101;
			10'b1101001011 		: log = 16'b0011100011001110;
			10'b1101001100 		: log = 16'b0011100011001111;
			10'b1101001101 		: log = 16'b0011100011010000;
			10'b1101001110 		: log = 16'b0011100011010001;
			10'b1101001111 		: log = 16'b0011100011010010;
			10'b1101010000 		: log = 16'b0011100011010100;
			10'b1101010001 		: log = 16'b0011100011010101;
			10'b1101010010 		: log = 16'b0011100011010110;
			10'b1101010011 		: log = 16'b0011100011010111;
			10'b1101010100 		: log = 16'b0011100011011000;
			10'b1101010101 		: log = 16'b0011100011011001;
			10'b1101010110 		: log = 16'b0011100011011010;
			10'b1101010111 		: log = 16'b0011100011011011;
			10'b1101011000 		: log = 16'b0011100011011100;
			10'b1101011001 		: log = 16'b0011100011011101;
			10'b1101011010 		: log = 16'b0011100011011110;
			10'b1101011011 		: log = 16'b0011100011100000;
			10'b1101011100 		: log = 16'b0011100011100001;
			10'b1101011101 		: log = 16'b0011100011100010;
			10'b1101011110 		: log = 16'b0011100011100011;
			10'b1101011111 		: log = 16'b0011100011100100;
			10'b1101100000 		: log = 16'b0011100011100101;
			10'b1101100001 		: log = 16'b0011100011100110;
			10'b1101100010 		: log = 16'b0011100011100111;
			10'b1101100011 		: log = 16'b0011100011101000;
			10'b1101100100 		: log = 16'b0011100011101001;
			10'b1101100101 		: log = 16'b0011100011101010;
			10'b1101100110 		: log = 16'b0011100011101011;
			10'b1101100111 		: log = 16'b0011100011101101;
			10'b1101101000 		: log = 16'b0011100011101110;
			10'b1101101001 		: log = 16'b0011100011101111;
			10'b1101101010 		: log = 16'b0011100011110000;
			10'b1101101011 		: log = 16'b0011100011110001;
			10'b1101101100 		: log = 16'b0011100011110010;
			10'b1101101101 		: log = 16'b0011100011110011;
			10'b1101101110 		: log = 16'b0011100011110100;
			10'b1101101111 		: log = 16'b0011100011110101;
			10'b1101110000 		: log = 16'b0011100011110110;
			10'b1101110001 		: log = 16'b0011100011110111;
			10'b1101110010 		: log = 16'b0011100011111000;
			10'b1101110011 		: log = 16'b0011100011111001;
			10'b1101110100 		: log = 16'b0011100011111011;
			10'b1101110101 		: log = 16'b0011100011111100;
			10'b1101110110 		: log = 16'b0011100011111101;
			10'b1101110111 		: log = 16'b0011100011111110;
			10'b1101111000 		: log = 16'b0011100011111111;
			10'b1101111001 		: log = 16'b0011100100000000;
			10'b1101111010 		: log = 16'b0011100100000001;
			10'b1101111011 		: log = 16'b0011100100000010;
			10'b1101111100 		: log = 16'b0011100100000011;
			10'b1101111101 		: log = 16'b0011100100000100;
			10'b1101111110 		: log = 16'b0011100100000101;
			10'b1101111111 		: log = 16'b0011100100000110;
			10'b1110000000 		: log = 16'b0011100100000111;
			10'b1110000001 		: log = 16'b0011100100001000;
			10'b1110000010 		: log = 16'b0011100100001010;
			10'b1110000011 		: log = 16'b0011100100001011;
			10'b1110000100 		: log = 16'b0011100100001100;
			10'b1110000101 		: log = 16'b0011100100001101;
			10'b1110000110 		: log = 16'b0011100100001110;
			10'b1110000111 		: log = 16'b0011100100001111;
			10'b1110001000 		: log = 16'b0011100100010000;
			10'b1110001001 		: log = 16'b0011100100010001;
			10'b1110001010 		: log = 16'b0011100100010010;
			10'b1110001011 		: log = 16'b0011100100010011;
			10'b1110001100 		: log = 16'b0011100100010100;
			10'b1110001101 		: log = 16'b0011100100010101;
			10'b1110001110 		: log = 16'b0011100100010110;
			10'b1110001111 		: log = 16'b0011100100010111;
			10'b1110010000 		: log = 16'b0011100100011000;
			10'b1110010001 		: log = 16'b0011100100011001;
			10'b1110010010 		: log = 16'b0011100100011011;
			10'b1110010011 		: log = 16'b0011100100011100;
			10'b1110010100 		: log = 16'b0011100100011101;
			10'b1110010101 		: log = 16'b0011100100011110;
			10'b1110010110 		: log = 16'b0011100100011111;
			10'b1110010111 		: log = 16'b0011100100100000;
			10'b1110011000 		: log = 16'b0011100100100001;
			10'b1110011001 		: log = 16'b0011100100100010;
			10'b1110011010 		: log = 16'b0011100100100011;
			10'b1110011011 		: log = 16'b0011100100100100;
			10'b1110011100 		: log = 16'b0011100100100101;
			10'b1110011101 		: log = 16'b0011100100100110;
			10'b1110011110 		: log = 16'b0011100100100111;
			10'b1110011111 		: log = 16'b0011100100101000;
			10'b1110100000 		: log = 16'b0011100100101001;
			10'b1110100001 		: log = 16'b0011100100101010;
			10'b1110100010 		: log = 16'b0011100100101011;
			10'b1110100011 		: log = 16'b0011100100101100;
			10'b1110100100 		: log = 16'b0011100100101101;
			10'b1110100101 		: log = 16'b0011100100101110;
			10'b1110100110 		: log = 16'b0011100100110000;
			10'b1110100111 		: log = 16'b0011100100110001;
			10'b1110101000 		: log = 16'b0011100100110010;
			10'b1110101001 		: log = 16'b0011100100110011;
			10'b1110101010 		: log = 16'b0011100100110100;
			10'b1110101011 		: log = 16'b0011100100110101;
			10'b1110101100 		: log = 16'b0011100100110110;
			10'b1110101101 		: log = 16'b0011100100110111;
			10'b1110101110 		: log = 16'b0011100100111000;
			10'b1110101111 		: log = 16'b0011100100111001;
			10'b1110110000 		: log = 16'b0011100100111010;
			10'b1110110001 		: log = 16'b0011100100111011;
			10'b1110110010 		: log = 16'b0011100100111100;
			10'b1110110011 		: log = 16'b0011100100111101;
			10'b1110110100 		: log = 16'b0011100100111110;
			10'b1110110101 		: log = 16'b0011100100111111;
			10'b1110110110 		: log = 16'b0011100101000000;
			10'b1110110111 		: log = 16'b0011100101000001;
			10'b1110111000 		: log = 16'b0011100101000010;
			10'b1110111001 		: log = 16'b0011100101000011;
			10'b1110111010 		: log = 16'b0011100101000100;
			10'b1110111011 		: log = 16'b0011100101000101;
			10'b1110111100 		: log = 16'b0011100101000110;
			10'b1110111101 		: log = 16'b0011100101000111;
			10'b1110111110 		: log = 16'b0011100101001000;
			10'b1110111111 		: log = 16'b0011100101001010;
			10'b1111000000 		: log = 16'b0011100101001011;
			10'b1111000001 		: log = 16'b0011100101001100;
			10'b1111000010 		: log = 16'b0011100101001101;
			10'b1111000011 		: log = 16'b0011100101001110;
			10'b1111000100 		: log = 16'b0011100101001111;
			10'b1111000101 		: log = 16'b0011100101010000;
			10'b1111000110 		: log = 16'b0011100101010001;
			10'b1111000111 		: log = 16'b0011100101010010;
			10'b1111001000 		: log = 16'b0011100101010011;
			10'b1111001001 		: log = 16'b0011100101010100;
			10'b1111001010 		: log = 16'b0011100101010101;
			10'b1111001011 		: log = 16'b0011100101010110;
			10'b1111001100 		: log = 16'b0011100101010111;
			10'b1111001101 		: log = 16'b0011100101011000;
			10'b1111001110 		: log = 16'b0011100101011001;
			10'b1111001111 		: log = 16'b0011100101011010;
			10'b1111010000 		: log = 16'b0011100101011011;
			10'b1111010001 		: log = 16'b0011100101011100;
			10'b1111010010 		: log = 16'b0011100101011101;
			10'b1111010011 		: log = 16'b0011100101011110;
			10'b1111010100 		: log = 16'b0011100101011111;
			10'b1111010101 		: log = 16'b0011100101100000;
			10'b1111010110 		: log = 16'b0011100101100001;
			10'b1111010111 		: log = 16'b0011100101100010;
			10'b1111011000 		: log = 16'b0011100101100011;
			10'b1111011001 		: log = 16'b0011100101100100;
			10'b1111011010 		: log = 16'b0011100101100101;
			10'b1111011011 		: log = 16'b0011100101100110;
			10'b1111011100 		: log = 16'b0011100101100111;
			10'b1111011101 		: log = 16'b0011100101101000;
			10'b1111011110 		: log = 16'b0011100101101001;
			10'b1111011111 		: log = 16'b0011100101101010;
			10'b1111100000 		: log = 16'b0011100101101011;
			10'b1111100001 		: log = 16'b0011100101101100;
			10'b1111100010 		: log = 16'b0011100101101101;
			10'b1111100011 		: log = 16'b0011100101101110;
			10'b1111100100 		: log = 16'b0011100101101111;
			10'b1111100101 		: log = 16'b0011100101110000;
			10'b1111100110 		: log = 16'b0011100101110001;
			10'b1111100111 		: log = 16'b0011100101110010;
			10'b1111101000 		: log = 16'b0011100101110011;
			10'b1111101001 		: log = 16'b0011100101110100;
			10'b1111101010 		: log = 16'b0011100101110101;
			10'b1111101011 		: log = 16'b0011100101110110;
			10'b1111101100 		: log = 16'b0011100101110111;
			10'b1111101101 		: log = 16'b0011100101111000;
			10'b1111101110 		: log = 16'b0011100101111001;
			10'b1111101111 		: log = 16'b0011100101111010;
			10'b1111110000 		: log = 16'b0011100101111100;
			10'b1111110001 		: log = 16'b0011100101111101;
			10'b1111110010 		: log = 16'b0011100101111110;
			10'b1111110011 		: log = 16'b0011100101111111;
			10'b1111110100 		: log = 16'b0011100110000000;
			10'b1111110101 		: log = 16'b0011100110000001;
			10'b1111110110 		: log = 16'b0011100110000010;
			10'b1111110111 		: log = 16'b0011100110000011;
			10'b1111111000 		: log = 16'b0011100110000100;
			10'b1111111001 		: log = 16'b0011100110000101;
			10'b1111111010 		: log = 16'b0011100110000110;
			10'b1111111011 		: log = 16'b0011100110000111;
			10'b1111111100 		: log = 16'b0011100110001000;
			10'b1111111101 		: log = 16'b0011100110001001;
			10'b1111111110 		: log = 16'b0011100110001010;
			10'b1111111111 		: log = 16'b0011100110001011;
        endcase
    end
endmodule
