`define DATAWIDTH 16

module mode2_sub(
  a_inp0,
  a_inp1,
  a_inp2,
  a_inp3,
  
  b_inp,
  
  outp0,
  outp1,
  outp2,
  outp3); 
  
  input  [`DATAWIDTH-1 : 0] a_inp0;
  input  [`DATAWIDTH-1 : 0] a_inp1;
  input  [`DATAWIDTH-1 : 0] a_inp2;
  input  [`DATAWIDTH-1 : 0] a_inp3;
  
  input  [`DATAWIDTH-1 : 0] b_inp;

  output [`DATAWIDTH-1 : 0] outp0;
  output [`DATAWIDTH-1 : 0] outp1;
  output [`DATAWIDTH-1 : 0] outp2;
  output [`DATAWIDTH-1 : 0] outp3;
  
  DW_fp_sub sub0(.a(a_inp0), .b(b_inp), .z(outp0), .rnd(3'b000));
  DW_fp_sub sub1(.a(a_inp1), .b(b_inp), .z(outp1), .rnd(3'b000));
  DW_fp_sub sub2(.a(a_inp2), .b(b_inp), .z(outp2), .rnd(3'b000));
  DW_fp_sub sub3(.a(a_inp3), .b(b_inp), .z(outp3), .rnd(3'b000));

endmodule

