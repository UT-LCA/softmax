module expunit (a, z, status, stage_run, clk, reset);

	parameter int_width = 3; // fixed point integer length
	parameter frac_width = 4; // fixed point fraction length
		
	input [31:0] a;
	input stage_run;
  	input clk;
  	input reset;
	output [31:0] z;
	output [7:0] status;
	//wire [int_width + frac_width - 1: 0] fxout;
	wire [63:0] LUTout;
	wire [63:0] Mult_out;
	reg [31:0] LUTout_reg;
	reg [31:0] Mult_out_reg;
	wire [int_width + frac_width - 1:0] fx;

	always @(posedge clk) begin
    		if(reset) begin
      		Mult_out_reg <= 0;
      		LUTout_reg <= 0;
    		end else if(stage_run) begin
      		Mult_out_reg <= Mult_out[47:16];
      		LUTout_reg <= LUTout[31:0];
    		end
  	end

	//fptofixed_para fpfx (.fp(a), .fx(fxout));
	fptofixed_para fptofx(.fp(a),.fx(fx));
	LUT lut(.addr(fx), .exp(LUTout)); 
	DW02_mult #(32,32) mult (.A(a), .B(LUTout[63:32]), .TC(1'b1), .PRODUCT(Mult_out));
	DW01_add #(32) add (.A(Mult_out_reg[31:0]), .B(LUTout_reg[31:0]), .CI(1'b0), .SUM(z), .CO());
endmodule

module fptofixed_para (
	fp,
	fx
	);
	
	parameter int_width = 3; // fixed point integer length
	parameter frac_width = 4; // fixed point fraction length

	input [31:0] fp; // Half Precision fp
	output [int_width + frac_width - 1:0] fx;  
	
	//wire [15:0] Mant; // mantissa of fp
	//wire signed [4:0] Ea; // non biased exponent
	//wire [4:0] Exp; // biased exponent
	//wire [15:0] sftfx; // output of shifter block
	wire [31:0] temp;
	wire grt;
	wire [31:0] temp2;
	reg [31:0] temp3;
	//assign Mant = {6'b000001, fp[9:0]};
	//assign Exp = fp[14:10];
	//assign Ea = Exp - 15;

	assign fx = temp3[15+int_width:16-frac_width];
	assign grt = |(temp2[31:16+int_width]);
	//assign neg = &(fp[31:16+int_width]);
	assign temp2 = ~(temp[31:0]);	

always @(temp2)
begin
// only negetive numbers as inputs after sorting and subtraction from max
	if (grt)
		begin
			temp3 <= 32'hFFFF; // if there is an overflow
			
		end
	//else if ( fp[14:0] == 15'b0)
	//	begin 
	//		temp <= 16'b0;
			
	
	else // underflow automatically becomes zero
		begin
			temp3 <= temp2;

		end
end	


//DW01_ash ash( .A(Mant[15:0]), .DATA_TC(1'b0), .SH(Ea[4:0]), .SH_TC(1'b1), .B(sftfx));
DW01_addsub #(32) addsub1 (.A(fp),.B(32'h00000001),.CI(1'b0),.ADD_SUB(1'b1),.SUM(temp),.CO());
endmodule

module LUT(addr, exp);
    input [6:0] addr;
    output reg [63:0] exp;

    always @(addr) begin
        case (addr)
	     7'b0000000            : exp =  64'b0000000000000000111110000010101000000000000000010000000000000000;
	     7'b0000001            : exp =  64'b0000000000000000111010010010000000000000000000001111111100001111;
	     7'b0000010            : exp =  64'b0000000000000000110110110000000100000000000000001111110101001011;
	     7'b0000011            : exp =  64'b0000000000000000110011011011110000000000000000001111101011001110;
	     7'b0000100            : exp =  64'b0000000000000000110000010100010100000000000000001111011110110000;
	     7'b0000101            : exp =  64'b0000000000000000101101011000111100000000000000001111010000001000;
	     7'b0000110            : exp =  64'b0000000000000000101010101000111100000000000000001110111111101000;
	     7'b0000111            : exp =  64'b0000000000000000101000000011101000000000000000001110101101100010;
	     7'b0001000            : exp =  64'b0000000000000000100101101000010000000000000000001110011010001000;
	     7'b0001001            : exp =  64'b0000000000000000100011010110011000000000000000001110000101100110;
	     7'b0001010            : exp =  64'b0000000000000000100001001101010100000000000000001101110000001100;
	     7'b0001011            : exp =  64'b0000000000000000011111001100100000000000000000001101011010000011;
	     7'b0001100            : exp =  64'b0000000000000000011101010011100100000000000000001101000011011000;
	     7'b0001101            : exp =  64'b0000000000000000011011100001111100000000000000001100101100010010;
	     7'b0001110            : exp =  64'b0000000000000000011001110111001100000000000000001100010100111100;
	     7'b0001111            : exp =  64'b0000000000000000011000010010111000000000000000001011111101011100;
	     7'b0010000            : exp =  64'b0000000000000000010110110100101100000000000000001011100101111000;
	     7'b0010001            : exp =  64'b0000000000000000010101011100001100000000000000001011001110011000;
	     7'b0010010            : exp =  64'b0000000000000000010100001001000100000000000000001010110110111111;
	     7'b0010011            : exp =  64'b0000000000000000010010111010111100000000000000001010011111110011;
	     7'b0010100            : exp =  64'b0000000000000000010001110001100100000000000000001010001000111000;
	     7'b0010101            : exp =  64'b0000000000000000010000101100101000000000000000001001110010010001;
	     7'b0010110            : exp =  64'b0000000000000000001111101011111000000000000000001001011100000000;
	     7'b0010111            : exp =  64'b0000000000000000001110101111000100000000000000001001000110001001;
	     7'b0011000            : exp =  64'b0000000000000000001101110101111100000000000000001000110000101110;
	     7'b0011001            : exp =  64'b0000000000000000001101000000010000000000000000001000011011110000;
	     7'b0011010            : exp =  64'b0000000000000000001100001101110100000000000000001000000111010001;
	     7'b0011011            : exp =  64'b0000000000000000001011011110011100000000000000000111110011010010;
	     7'b0011100            : exp =  64'b0000000000000000001010110001111100000000000000000111011111110100;
	     7'b0011101            : exp =  64'b0000000000000000001010001000001000000000000000000111001100110111;
	     7'b0011110            : exp =  64'b0000000000000000001001100000111000000000000000000110111010011101;
	     7'b0011111            : exp =  64'b0000000000000000001000111100000000000000000000000110101000100110;
	     7'b0100000            : exp =  64'b0000000000000000001000011001010100000000000000000110010111010001;
	     7'b0100001            : exp =  64'b0000000000000000000111111000110000000000000000000110000110011110;
	     7'b0100010            : exp =  64'b0000000000000000000111011010001100000000000000000101110110001110;
	     7'b0100011            : exp =  64'b0000000000000000000110111101011100000000000000000101100110100001;
	     7'b0100100            : exp =  64'b0000000000000000000110100010100000000000000000000101010111010101;
	     7'b0100101            : exp =  64'b0000000000000000000110001001001000000000000000000101001000101011;
	     7'b0100110            : exp =  64'b0000000000000000000101110001010100000000000000000100111010100010;
	     7'b0100111            : exp =  64'b0000000000000000000101011010111100000000000000000100101100111001;
	     7'b0101000            : exp =  64'b0000000000000000000101000101111000000000000000000100011111110000;
	     7'b0101001            : exp =  64'b0000000000000000000100110010001000000000000000000100010011000111;
	     7'b0101010            : exp =  64'b0000000000000000000100011111101000000000000000000100000110111011;
	     7'b0101011            : exp =  64'b0000000000000000000100001110001100000000000000000011111011001110;
	     7'b0101100            : exp =  64'b0000000000000000000011111101110100000000000000000011101111111110;
	     7'b0101101            : exp =  64'b0000000000000000000011101110011100000000000000000011100101001010;
	     7'b0101110            : exp =  64'b0000000000000000000011100000000000000000000000000011011010110001;
	     7'b0101111            : exp =  64'b0000000000000000000011010010011000000000000000000011010000110011;
	     7'b0110000            : exp =  64'b0000000000000000000011000101101000000000000000000011000111001111;
	     7'b0110001            : exp =  64'b0000000000000000000010111001101100000000000000000010111110000100;
	     7'b0110010            : exp =  64'b0000000000000000000010101110011100000000000000000010110101010010;
	     7'b0110011            : exp =  64'b0000000000000000000010100011111000000000000000000010101100110111;
	     7'b0110100            : exp =  64'b0000000000000000000010011001111100000000000000000010100100110010;
	     7'b0110101            : exp =  64'b0000000000000000000010010000101000000000000000000010011101000100;
	     7'b0110110            : exp =  64'b0000000000000000000010000111110100000000000000000010010101101011;
	     7'b0110111            : exp =  64'b0000000000000000000001111111101000000000000000000010001110100110;
	     7'b0111000            : exp =  64'b0000000000000000000001110111111000000000000000000010000111110101;
	     7'b0111001            : exp =  64'b0000000000000000000001110000101000000000000000000010000001010111;
	     7'b0111010            : exp =  64'b0000000000000000000001101001110100000000000000000001111011001011;
	     7'b0111011            : exp =  64'b0000000000000000000001100011011000000000000000000001110101010001;
	     7'b0111100            : exp =  64'b0000000000000000000001011101011000000000000000000001101111101000;
	     7'b0111101            : exp =  64'b0000000000000000000001010111101100000000000000000001101010001110;
	     7'b0111110            : exp =  64'b0000000000000000000001010010011000000000000000000001100101000101;
	     7'b0111111            : exp =  64'b0000000000000000000001001101011000000000000000000001100000001010;
	     7'b1000000            : exp =  64'b0000000000000000000001001000101100000000000000000001011011011110;
	     7'b1000001            : exp =  64'b0000000000000000000001000100010100000000000000000001010111000000;
	     7'b1000010            : exp =  64'b0000000000000000000001000000001000000000000000000001010010101111;
	     7'b1000011            : exp =  64'b0000000000000000000000111100010000000000000000000001001110101010;
	     7'b1000100            : exp =  64'b0000000000000000000000111000101000000000000000000001001010110010;
	     7'b1000101            : exp =  64'b0000000000000000000000110101001100000000000000000001000111000101;
	     7'b1000110            : exp =  64'b0000000000000000000000110001111100000000000000000001000011100011;
	     7'b1000111            : exp =  64'b0000000000000000000000101110111100000000000000000001000000001100;
	     7'b1001000            : exp =  64'b0000000000000000000000101100000100000000000000000000111100111111;
	     7'b1001001            : exp =  64'b0000000000000000000000101001011000000000000000000000111001111100;
	     7'b1001010            : exp =  64'b0000000000000000000000100110111000000000000000000000110111000011;
	     7'b1001011            : exp =  64'b0000000000000000000000100100100100000000000000000000110100010010;
	     7'b1001100            : exp =  64'b0000000000000000000000100010010100000000000000000000110001101001;
	     7'b1001101            : exp =  64'b0000000000000000000000100000010000000000000000000000101111001001;
	     7'b1001110            : exp =  64'b0000000000000000000000011110010100000000000000000000101100110001;
	     7'b1001111            : exp =  64'b0000000000000000000000011100011100000000000000000000101010011111;
	     7'b1010000            : exp =  64'b0000000000000000000000011010110000000000000000000000101000010101;
	     7'b1010001            : exp =  64'b0000000000000000000000011001001000000000000000000000100110010010;
	     7'b1010010            : exp =  64'b0000000000000000000000010111100100000000000000000000100100010101;
	     7'b1010011            : exp =  64'b0000000000000000000000010110001000000000000000000000100010011110;
	     7'b1010100            : exp =  64'b0000000000000000000000010100110100000000000000000000100000101110;
	     7'b1010101            : exp =  64'b0000000000000000000000010011100100000000000000000000011111000010;
	     7'b1010110            : exp =  64'b0000000000000000000000010010011000000000000000000000011101011100;
	     7'b1010111            : exp =  64'b0000000000000000000000010001010000000000000000000000011011111011;
	     7'b1011000            : exp =  64'b0000000000000000000000010000001100000000000000000000011010011111;
	     7'b1011001            : exp =  64'b0000000000000000000000001111001100000000000000000000011001001000;
	     7'b1011010            : exp =  64'b0000000000000000000000001110010100000000000000000000010111110101;
	     7'b1011011            : exp =  64'b0000000000000000000000001101011100000000000000000000010110100110;
	     7'b1011100            : exp =  64'b0000000000000000000000001100101000000000000000000000010101011011;
	     7'b1011101            : exp =  64'b0000000000000000000000001011110100000000000000000000010100010100;
	     7'b1011110            : exp =  64'b0000000000000000000000001011001000000000000000000000010011010000;
	     7'b1011111            : exp =  64'b0000000000000000000000001010011100000000000000000000010010010000;
	     7'b1100000            : exp =  64'b0000000000000000000000001001110100000000000000000000010001010011;
	     7'b1100001            : exp =  64'b0000000000000000000000001001001100000000000000000000010000011001;
	     7'b1100010            : exp =  64'b0000000000000000000000001000101000000000000000000000001111100010;
	     7'b1100011            : exp =  64'b0000000000000000000000001000001000000000000000000000001110101110;
	     7'b1100100            : exp =  64'b0000000000000000000000000111101000000000000000000000001101111101;
	     7'b1100101            : exp =  64'b0000000000000000000000000111001100000000000000000000001101001110;
	     7'b1100110            : exp =  64'b0000000000000000000000000110110000000000000000000000001100100001;
	     7'b1100111            : exp =  64'b0000000000000000000000000110010100000000000000000000001011110111;
	     7'b1101000            : exp =  64'b0000000000000000000000000101111100000000000000000000001011001111;
	     7'b1101001            : exp =  64'b0000000000000000000000000101100100000000000000000000001010101001;
	     7'b1101010            : exp =  64'b0000000000000000000000000101010000000000000000000000001010000101;
	     7'b1101011            : exp =  64'b0000000000000000000000000100111100000000000000000000001001100011;
	     7'b1101100            : exp =  64'b0000000000000000000000000100101000000000000000000000001001000010;
	     7'b1101101            : exp =  64'b0000000000000000000000000100010100000000000000000000001000100100;
	     7'b1101110            : exp =  64'b0000000000000000000000000100000100000000000000000000001000000111;
	     7'b1101111            : exp =  64'b0000000000000000000000000011110100000000000000000000000111101011;
	     7'b1110000            : exp =  64'b0000000000000000000000000011100100000000000000000000000111010001;
	     7'b1110001            : exp =  64'b0000000000000000000000000011011000000000000000000000000110111000;
	     7'b1110010            : exp =  64'b0000000000000000000000000011001100000000000000000000000110100001;
	     7'b1110011            : exp =  64'b0000000000000000000000000011000000000000000000000000000110001010;
	     7'b1110100            : exp =  64'b0000000000000000000000000010110100000000000000000000000101110101;
	     7'b1110101            : exp =  64'b0000000000000000000000000010101000000000000000000000000101100001;
	     7'b1110110            : exp =  64'b0000000000000000000000000010011100000000000000000000000101001110;
	     7'b1110111            : exp =  64'b0000000000000000000000000010010100000000000000000000000100111100;
	     7'b1111000            : exp =  64'b0000000000000000000000000010001100000000000000000000000100101011;
	     7'b1111001            : exp =  64'b0000000000000000000000000010000100000000000000000000000100011011;
	     7'b1111010            : exp =  64'b0000000000000000000000000001111100000000000000000000000100001100;
	     7'b1111011            : exp =  64'b0000000000000000000000000001110100000000000000000000000011111101;
	     7'b1111100            : exp =  64'b0000000000000000000000000001101100000000000000000000000011110000;
	     7'b1111101            : exp =  64'b0000000000000000000000000001100100000000000000000000000011100011;
	     7'b1111110            : exp =  64'b0000000000000000000000000001100000000000000000000000000011010111;
	     7'b1111111            : exp =  64'b0000000000000000000000000001011000000000000000000000000011001011;
        endcase
    end
endmodule
