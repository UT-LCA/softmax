module LUT2(addr, log);
    input [5:0] addr;
    output reg [15:0] log;

    always @(addr) begin
        case (addr)
			5'b0 		: log = 16'b0000000000000000;
			5'b1 		: log = 16'b0010001111110000;
			5'b10 		: log = 16'b0010011111100001;
			5'b11 		: log = 16'b0010100111011101;
			5'b100 		: log = 16'b0010101111000011;
			5'b101 		: log = 16'b0010110011010000;
			5'b110 		: log = 16'b0010110110111100;
			5'b111 		: log = 16'b0010111010100101;
			5'b1000 		: log = 16'b0010111110001010;
			5'b1001 		: log = 16'b0011000000110110;
			5'b1010 		: log = 16'b0011000010100101;
			5'b1011 		: log = 16'b0011000100010011;
			5'b1100 		: log = 16'b0011000110000000;
			5'b1101 		: log = 16'b0011000111101011;
			5'b1110 		: log = 16'b0011001001010101;
			5'b1111 		: log = 16'b0011001010111101;
			5'b10000 		: log = 16'b0011001100100100;
			5'b10001 		: log = 16'b0011001110001010;
			5'b10010 		: log = 16'b0011001111101110;
			5'b10011 		: log = 16'b0011010000101001;
			5'b10100 		: log = 16'b0011010001011010;
			5'b10101 		: log = 16'b0011010010001010;
			5'b10110 		: log = 16'b0011010010111010;
			5'b10111 		: log = 16'b0011010011101010;
			5'b11000 		: log = 16'b0011010100011000;
			5'b11001 		: log = 16'b0011010101000111;
			5'b11010 		: log = 16'b0011010101110100;
			5'b11011 		: log = 16'b0011010110100010;
			5'b11100 		: log = 16'b0011010111001110;
			5'b11101 		: log = 16'b0011010111111011;
			5'b11110 		: log = 16'b0011011000100111;
			5'b11111 		: log = 16'b0011011001010010;
			5'b100000 		: log = 16'b0011011001111101;
			5'b100001 		: log = 16'b0011011010100111;
			5'b100010 		: log = 16'b0011011011010001;
			5'b100011 		: log = 16'b0011011011111011;
			5'b100100 		: log = 16'b0011011100100100;
			5'b100101 		: log = 16'b0011011101001101;
			5'b100110 		: log = 16'b0011011101110101;
			5'b100111 		: log = 16'b0011011110011101;
			5'b101000 		: log = 16'b0011011111000101;
			5'b101001 		: log = 16'b0011011111101100;
			5'b101010 		: log = 16'b0011100000001001;
			5'b101011 		: log = 16'b0011100000011101;
			5'b101100 		: log = 16'b0011100000110000;
			5'b101101 		: log = 16'b0011100001000010;
			5'b101110 		: log = 16'b0011100001010101;
			5'b101111 		: log = 16'b0011100001101000;
			5'b110000 		: log = 16'b0011100001111010;
			5'b110001 		: log = 16'b0011100010001100;
			5'b110010 		: log = 16'b0011100010011110;
			5'b110011 		: log = 16'b0011100010110000;
			5'b110100 		: log = 16'b0011100011000010;
			5'b110101 		: log = 16'b0011100011010100;
			5'b110110 		: log = 16'b0011100011100101;
			5'b110111 		: log = 16'b0011100011110110;
			5'b111000 		: log = 16'b0011100100000111;
			5'b111001 		: log = 16'b0011100100011000;
			5'b111010 		: log = 16'b0011100100101001;
			5'b111011 		: log = 16'b0011100100111010;
			5'b111100 		: log = 16'b0011100101001011;
			5'b111101 		: log = 16'b0011100101011011;
			5'b111110 		: log = 16'b0011100101101011;
			5'b111111 		: log = 16'b0011100101111100;
        endcase
    end
endmodule
